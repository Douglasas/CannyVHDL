library ieee;
use ieee.std_logic_1164.all;

package main_pkg is
  constant INPUT_IMAGE_X : integer := 481;
  constant INPUT_IMAGE_Y : integer := 321;
end package;
