library ieee;
use ieee.std_logic_1164.all;

package main_pkg is
  constant INPUT_IMAGE_Y : integer := 512;
  constant INPUT_IMAGE_X : integer := 512;
end package;
