-- megafunction wizard: %ALTSQRT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTSQRT

-- ============================================================
-- File Name: sqrtip.vhd
-- Megafunction Name(s):
-- 			ALTSQRT
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.4 Build 182 03/12/2014 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2014 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions
--and other software and tools, and its AMPP partner logic
--functions, and any output files from any of the foregoing
--(including device programming or simulation files), and any
--associated documentation or information are expressly subject
--to the terms and conditions of the Altera Program License
--Subscription Agreement, Altera MegaCore Function License
--Agreement, or other applicable license agreement, including,
--without limitation, that your use is for the sole purpose of
--programming logic devices manufactured by Altera and sold by
--Altera or its authorized distributors.  Please refer to the
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

library work;
use work.slogic_pkg.all;
use work.gradient_pkg.all;

ENTITY sqrtip IS
	PORT
	(
		clk		: IN STD_LOGIC ;
		ena		: IN STD_LOGIC ;
		radical		: IN STD_LOGIC_VECTOR (2*(MSB+LSB)-1 DOWNTO 0);
		q		: OUT STD_LOGIC_VECTOR (MSB+LSB-1 DOWNTO 0);
		remainder		: OUT STD_LOGIC_VECTOR (MSB+LSB DOWNTO 0)
	);
END sqrtip;


ARCHITECTURE SYN OF sqrtip IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (MSB+LSB-1 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (MSB+LSB DOWNTO 0);



	COMPONENT altsqrt
	GENERIC (
		pipeline     : NATURAL;
		q_port_width : NATURAL;
		r_port_width : NATURAL;
		width        : NATURAL;
		lpm_type		 : STRING
	);
	PORT (
			clk	: IN STD_LOGIC ;
			ena	: IN STD_LOGIC ;
			radical	: IN STD_LOGIC_VECTOR (2*(MSB+LSB)-1 DOWNTO 0);
			q	: OUT STD_LOGIC_VECTOR (MSB+LSB-1 DOWNTO 0);
			remainder	: OUT STD_LOGIC_VECTOR (MSB+LSB DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	q    <= sub_wire0(MSB+LSB-1 DOWNTO 0);
	remainder    <= sub_wire1(MSB+LSB DOWNTO 0);

	ALTSQRT_component : ALTSQRT
	GENERIC MAP (
		pipeline => QT_SQRT_CYCLES,
		q_port_width => MSB+LSB,
		r_port_width => MSB+LSB+1,
		width => 2*(MSB+LSB),
		lpm_type => "ALTSQRT"
	)
	PORT MAP (
		clk => clk,
		ena => ena,
		radical => radical,
		q => sub_wire0,
		remainder => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "10"
-- Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "34"
-- Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "35"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "68"
-- Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL "clk"
-- Retrieval info: USED_PORT: ena 0 0 0 0 INPUT NODEFVAL "ena"
-- Retrieval info: USED_PORT: q 0 0 34 0 OUTPUT NODEFVAL "q[33..0]"
-- Retrieval info: USED_PORT: radical 0 0 68 0 INPUT NODEFVAL "radical[67..0]"
-- Retrieval info: USED_PORT: remainder 0 0 35 0 OUTPUT NODEFVAL "remainder[34..0]"
-- Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
-- Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
-- Retrieval info: CONNECT: @radical 0 0 68 0 radical 0 0 68 0
-- Retrieval info: CONNECT: q 0 0 34 0 @q 0 0 34 0
-- Retrieval info: CONNECT: remainder 0 0 35 0 @remainder 0 0 35 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL sqrtip.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sqrtip.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sqrtip.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sqrtip.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sqrtip_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
