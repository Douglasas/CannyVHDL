library ieee;
use ieee.std_logic_1164.all;

package main_pkg is
  constant INPUT_IMAGE_X : integer := 220;
  constant INPUT_IMAGE_Y : integer := 220;
end package;
