library ieee;
use ieee.std_logic_1164;
use ieee.numeric_std.all;

library work;
use work.main_pkg.all;
use work.slogic_pkg.all;

package tests_pkg is

  constant IMAGE_DATA : slogic_vec (0 to INPUT_IMAGE_X*INPUT_IMAGE_Y-1) := (
    to_slogic(157),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(150),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(144),
    to_slogic(146),
    to_slogic(126),
    to_slogic(102),
    to_slogic(87),
    to_slogic(96),
    to_slogic(96),
    to_slogic(109),
    to_slogic(103),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(121),
    to_slogic(118),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(135),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(130),
    to_slogic(139),
    to_slogic(128),
    to_slogic(135),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(128),
    to_slogic(135),
    to_slogic(130),
    to_slogic(126),
    to_slogic(133),
    to_slogic(133),
    to_slogic(134),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(135),
    to_slogic(126),
    to_slogic(133),
    to_slogic(137),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(128),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(133),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(107),
    to_slogic(109),
    to_slogic(101),
    to_slogic(116),
    to_slogic(126),
    to_slogic(144),
    to_slogic(137),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(158),
    to_slogic(158),
    to_slogic(157),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(150),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(156),
    to_slogic(152),
    to_slogic(156),
    to_slogic(144),
    to_slogic(157),
    to_slogic(144),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(158),
    to_slogic(157),
    to_slogic(156),
    to_slogic(150),
    to_slogic(178),
    to_slogic(205),
    to_slogic(207),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(197),
    to_slogic(150),
    to_slogic(101),
    to_slogic(101),
    to_slogic(109),
    to_slogic(107),
    to_slogic(118),
    to_slogic(117),
    to_slogic(128),
    to_slogic(124),
    to_slogic(117),
    to_slogic(126),
    to_slogic(118),
    to_slogic(128),
    to_slogic(118),
    to_slogic(117),
    to_slogic(126),
    to_slogic(117),
    to_slogic(124),
    to_slogic(118),
    to_slogic(126),
    to_slogic(126),
    to_slogic(118),
    to_slogic(128),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(118),
    to_slogic(128),
    to_slogic(126),
    to_slogic(118),
    to_slogic(126),
    to_slogic(118),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(133),
    to_slogic(162),
    to_slogic(173),
    to_slogic(144),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(165),
    to_slogic(172),
    to_slogic(157),
    to_slogic(152),
    to_slogic(146),
    to_slogic(117),
    to_slogic(102),
    to_slogic(102),
    to_slogic(81),
    to_slogic(102),
    to_slogic(103),
    to_slogic(101),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(116),
    to_slogic(117),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(121),
    to_slogic(133),
    to_slogic(130),
    to_slogic(134),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(135),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(130),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(130),
    to_slogic(128),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(139),
    to_slogic(130),
    to_slogic(133),
    to_slogic(134),
    to_slogic(133),
    to_slogic(144),
    to_slogic(130),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(133),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(118),
    to_slogic(119),
    to_slogic(119),
    to_slogic(126),
    to_slogic(117),
    to_slogic(107),
    to_slogic(109),
    to_slogic(100),
    to_slogic(117),
    to_slogic(118),
    to_slogic(139),
    to_slogic(137),
    to_slogic(152),
    to_slogic(150),
    to_slogic(165),
    to_slogic(157),
    to_slogic(158),
    to_slogic(157),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(150),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(150),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(184),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(197),
    to_slogic(150),
    to_slogic(107),
    to_slogic(102),
    to_slogic(101),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(118),
    to_slogic(128),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(117),
    to_slogic(118),
    to_slogic(124),
    to_slogic(118),
    to_slogic(128),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(118),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(162),
    to_slogic(173),
    to_slogic(144),
    to_slogic(165),
    to_slogic(155),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(151),
    to_slogic(156),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(139),
    to_slogic(118),
    to_slogic(102),
    to_slogic(87),
    to_slogic(103),
    to_slogic(92),
    to_slogic(96),
    to_slogic(102),
    to_slogic(101),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(135),
    to_slogic(135),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(128),
    to_slogic(135),
    to_slogic(128),
    to_slogic(135),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(135),
    to_slogic(126),
    to_slogic(130),
    to_slogic(137),
    to_slogic(128),
    to_slogic(126),
    to_slogic(135),
    to_slogic(126),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(128),
    to_slogic(133),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(118),
    to_slogic(119),
    to_slogic(107),
    to_slogic(116),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(126),
    to_slogic(130),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(155),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(156),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(156),
    to_slogic(157),
    to_slogic(151),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(144),
    to_slogic(150),
    to_slogic(172),
    to_slogic(197),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(222),
    to_slogic(205),
    to_slogic(172),
    to_slogic(118),
    to_slogic(101),
    to_slogic(109),
    to_slogic(107),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(126),
    to_slogic(118),
    to_slogic(128),
    to_slogic(118),
    to_slogic(117),
    to_slogic(126),
    to_slogic(118),
    to_slogic(117),
    to_slogic(128),
    to_slogic(126),
    to_slogic(118),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(128),
    to_slogic(118),
    to_slogic(126),
    to_slogic(126),
    to_slogic(118),
    to_slogic(126),
    to_slogic(118),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(124),
    to_slogic(137),
    to_slogic(128),
    to_slogic(83),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(152),
    to_slogic(156),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(144),
    to_slogic(135),
    to_slogic(117),
    to_slogic(102),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(107),
    to_slogic(116),
    to_slogic(116),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(135),
    to_slogic(133),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(130),
    to_slogic(133),
    to_slogic(134),
    to_slogic(130),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(135),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(134),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(128),
    to_slogic(117),
    to_slogic(117),
    to_slogic(107),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(128),
    to_slogic(133),
    to_slogic(137),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(151),
    to_slogic(144),
    to_slogic(156),
    to_slogic(152),
    to_slogic(156),
    to_slogic(144),
    to_slogic(157),
    to_slogic(151),
    to_slogic(156),
    to_slogic(150),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(156),
    to_slogic(183),
    to_slogic(203),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(191),
    to_slogic(143),
    to_slogic(109),
    to_slogic(101),
    to_slogic(117),
    to_slogic(107),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(117),
    to_slogic(118),
    to_slogic(128),
    to_slogic(117),
    to_slogic(128),
    to_slogic(119),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(118),
    to_slogic(126),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(109),
    to_slogic(75),
    to_slogic(56),
    to_slogic(49),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(156),
    to_slogic(151),
    to_slogic(165),
    to_slogic(161),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(169),
    to_slogic(165),
    to_slogic(151),
    to_slogic(144),
    to_slogic(130),
    to_slogic(117),
    to_slogic(102),
    to_slogic(92),
    to_slogic(81),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(94),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(135),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(133),
    to_slogic(135),
    to_slogic(126),
    to_slogic(135),
    to_slogic(133),
    to_slogic(134),
    to_slogic(130),
    to_slogic(139),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(128),
    to_slogic(130),
    to_slogic(133),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(128),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(119),
    to_slogic(133),
    to_slogic(139),
    to_slogic(151),
    to_slogic(152),
    to_slogic(155),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(157),
    to_slogic(156),
    to_slogic(151),
    to_slogic(157),
    to_slogic(156),
    to_slogic(143),
    to_slogic(156),
    to_slogic(157),
    to_slogic(152),
    to_slogic(156),
    to_slogic(156),
    to_slogic(152),
    to_slogic(158),
    to_slogic(191),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(205),
    to_slogic(184),
    to_slogic(118),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(107),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(126),
    to_slogic(119),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(118),
    to_slogic(126),
    to_slogic(118),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(118),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(118),
    to_slogic(101),
    to_slogic(75),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(165),
    to_slogic(158),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(161),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(143),
    to_slogic(135),
    to_slogic(116),
    to_slogic(102),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(130),
    to_slogic(134),
    to_slogic(126),
    to_slogic(133),
    to_slogic(128),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(126),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(134),
    to_slogic(128),
    to_slogic(135),
    to_slogic(128),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(135),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(126),
    to_slogic(135),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(117),
    to_slogic(126),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(101),
    to_slogic(101),
    to_slogic(117),
    to_slogic(128),
    to_slogic(137),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(156),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(144),
    to_slogic(156),
    to_slogic(143),
    to_slogic(144),
    to_slogic(157),
    to_slogic(176),
    to_slogic(197),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(197),
    to_slogic(158),
    to_slogic(107),
    to_slogic(109),
    to_slogic(107),
    to_slogic(117),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(117),
    to_slogic(117),
    to_slogic(126),
    to_slogic(128),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(109),
    to_slogic(75),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(158),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(157),
    to_slogic(156),
    to_slogic(143),
    to_slogic(130),
    to_slogic(117),
    to_slogic(102),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(96),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(116),
    to_slogic(128),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(134),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(133),
    to_slogic(128),
    to_slogic(133),
    to_slogic(130),
    to_slogic(126),
    to_slogic(128),
    to_slogic(134),
    to_slogic(133),
    to_slogic(128),
    to_slogic(135),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(130),
    to_slogic(135),
    to_slogic(133),
    to_slogic(139),
    to_slogic(126),
    to_slogic(128),
    to_slogic(135),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(133),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(128),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(110),
    to_slogic(109),
    to_slogic(109),
    to_slogic(119),
    to_slogic(133),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(165),
    to_slogic(155),
    to_slogic(165),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(151),
    to_slogic(157),
    to_slogic(156),
    to_slogic(156),
    to_slogic(144),
    to_slogic(152),
    to_slogic(156),
    to_slogic(143),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(191),
    to_slogic(205),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(183),
    to_slogic(137),
    to_slogic(101),
    to_slogic(109),
    to_slogic(107),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(126),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(128),
    to_slogic(126),
    to_slogic(117),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(118),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(96),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(152),
    to_slogic(143),
    to_slogic(130),
    to_slogic(116),
    to_slogic(102),
    to_slogic(92),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(134),
    to_slogic(126),
    to_slogic(130),
    to_slogic(135),
    to_slogic(133),
    to_slogic(135),
    to_slogic(126),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(135),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(135),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(139),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(135),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(128),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(101),
    to_slogic(101),
    to_slogic(102),
    to_slogic(119),
    to_slogic(128),
    to_slogic(139),
    to_slogic(144),
    to_slogic(151),
    to_slogic(157),
    to_slogic(155),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(156),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(144),
    to_slogic(151),
    to_slogic(152),
    to_slogic(144),
    to_slogic(172),
    to_slogic(197),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(205),
    to_slogic(172),
    to_slogic(118),
    to_slogic(101),
    to_slogic(101),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(118),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(128),
    to_slogic(118),
    to_slogic(119),
    to_slogic(118),
    to_slogic(128),
    to_slogic(126),
    to_slogic(118),
    to_slogic(133),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(135),
    to_slogic(119),
    to_slogic(94),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(144),
    to_slogic(137),
    to_slogic(128),
    to_slogic(101),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(99),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(135),
    to_slogic(126),
    to_slogic(135),
    to_slogic(128),
    to_slogic(135),
    to_slogic(133),
    to_slogic(130),
    to_slogic(134),
    to_slogic(133),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(130),
    to_slogic(134),
    to_slogic(135),
    to_slogic(134),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(135),
    to_slogic(126),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(126),
    to_slogic(134),
    to_slogic(128),
    to_slogic(126),
    to_slogic(133),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(135),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(134),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(130),
    to_slogic(137),
    to_slogic(135),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(134),
    to_slogic(124),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(134),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(117),
    to_slogic(117),
    to_slogic(110),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(117),
    to_slogic(119),
    to_slogic(137),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(162),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(150),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(143),
    to_slogic(157),
    to_slogic(151),
    to_slogic(144),
    to_slogic(156),
    to_slogic(184),
    to_slogic(205),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(191),
    to_slogic(143),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(117),
    to_slogic(107),
    to_slogic(117),
    to_slogic(117),
    to_slogic(126),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(126),
    to_slogic(118),
    to_slogic(128),
    to_slogic(126),
    to_slogic(118),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(135),
    to_slogic(133),
    to_slogic(126),
    to_slogic(94),
    to_slogic(64),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(151),
    to_slogic(144),
    to_slogic(135),
    to_slogic(117),
    to_slogic(109),
    to_slogic(92),
    to_slogic(83),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(107),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(117),
    to_slogic(118),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(128),
    to_slogic(135),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(135),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(139),
    to_slogic(137),
    to_slogic(133),
    to_slogic(130),
    to_slogic(128),
    to_slogic(135),
    to_slogic(128),
    to_slogic(133),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(128),
    to_slogic(119),
    to_slogic(128),
    to_slogic(117),
    to_slogic(116),
    to_slogic(101),
    to_slogic(117),
    to_slogic(101),
    to_slogic(102),
    to_slogic(110),
    to_slogic(117),
    to_slogic(139),
    to_slogic(144),
    to_slogic(152),
    to_slogic(155),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(158),
    to_slogic(157),
    to_slogic(165),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(156),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(156),
    to_slogic(143),
    to_slogic(151),
    to_slogic(152),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(165),
    to_slogic(191),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(176),
    to_slogic(118),
    to_slogic(109),
    to_slogic(102),
    to_slogic(117),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(128),
    to_slogic(118),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(130),
    to_slogic(92),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(156),
    to_slogic(165),
    to_slogic(157),
    to_slogic(156),
    to_slogic(144),
    to_slogic(135),
    to_slogic(117),
    to_slogic(100),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(97),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(126),
    to_slogic(121),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(135),
    to_slogic(133),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(133),
    to_slogic(134),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(128),
    to_slogic(134),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(135),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(135),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(117),
    to_slogic(128),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(107),
    to_slogic(119),
    to_slogic(128),
    to_slogic(139),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(155),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(158),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(144),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(184),
    to_slogic(205),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(197),
    to_slogic(161),
    to_slogic(107),
    to_slogic(109),
    to_slogic(107),
    to_slogic(107),
    to_slogic(117),
    to_slogic(118),
    to_slogic(126),
    to_slogic(117),
    to_slogic(116),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(118),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(128),
    to_slogic(92),
    to_slogic(63),
    to_slogic(63),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(143),
    to_slogic(135),
    to_slogic(116),
    to_slogic(97),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(94),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(128),
    to_slogic(134),
    to_slogic(126),
    to_slogic(130),
    to_slogic(135),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(134),
    to_slogic(126),
    to_slogic(121),
    to_slogic(130),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(135),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(134),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(119),
    to_slogic(119),
    to_slogic(126),
    to_slogic(128),
    to_slogic(119),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(101),
    to_slogic(119),
    to_slogic(119),
    to_slogic(128),
    to_slogic(146),
    to_slogic(146),
    to_slogic(152),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(161),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(158),
    to_slogic(191),
    to_slogic(207),
    to_slogic(213),
    to_slogic(222),
    to_slogic(222),
    to_slogic(222),
    to_slogic(205),
    to_slogic(191),
    to_slogic(124),
    to_slogic(101),
    to_slogic(109),
    to_slogic(116),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(126),
    to_slogic(128),
    to_slogic(118),
    to_slogic(126),
    to_slogic(117),
    to_slogic(128),
    to_slogic(117),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(126),
    to_slogic(133),
    to_slogic(133),
    to_slogic(126),
    to_slogic(92),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(161),
    to_slogic(165),
    to_slogic(156),
    to_slogic(143),
    to_slogic(135),
    to_slogic(116),
    to_slogic(100),
    to_slogic(89),
    to_slogic(89),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(117),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(133),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(128),
    to_slogic(134),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(139),
    to_slogic(133),
    to_slogic(133),
    to_slogic(134),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(117),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(121),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(128),
    to_slogic(133),
    to_slogic(130),
    to_slogic(133),
    to_slogic(133),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(119),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(128),
    to_slogic(128),
    to_slogic(137),
    to_slogic(146),
    to_slogic(155),
    to_slogic(151),
    to_slogic(157),
    to_slogic(162),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(155),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(161),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(150),
    to_slogic(157),
    to_slogic(143),
    to_slogic(157),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(176),
    to_slogic(203),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(222),
    to_slogic(222),
    to_slogic(205),
    to_slogic(172),
    to_slogic(116),
    to_slogic(109),
    to_slogic(107),
    to_slogic(117),
    to_slogic(116),
    to_slogic(117),
    to_slogic(118),
    to_slogic(126),
    to_slogic(117),
    to_slogic(118),
    to_slogic(126),
    to_slogic(117),
    to_slogic(118),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(133),
    to_slogic(139),
    to_slogic(126),
    to_slogic(99),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(156),
    to_slogic(143),
    to_slogic(135),
    to_slogic(121),
    to_slogic(94),
    to_slogic(92),
    to_slogic(82),
    to_slogic(99),
    to_slogic(96),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(124),
    to_slogic(118),
    to_slogic(121),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(134),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(134),
    to_slogic(135),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(133),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(133),
    to_slogic(128),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(121),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(110),
    to_slogic(110),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(155),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(152),
    to_slogic(150),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(157),
    to_slogic(191),
    to_slogic(203),
    to_slogic(203),
    to_slogic(222),
    to_slogic(222),
    to_slogic(222),
    to_slogic(213),
    to_slogic(197),
    to_slogic(143),
    to_slogic(110),
    to_slogic(110),
    to_slogic(110),
    to_slogic(116),
    to_slogic(116),
    to_slogic(117),
    to_slogic(118),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(118),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(130),
    to_slogic(133),
    to_slogic(118),
    to_slogic(92),
    to_slogic(50),
    to_slogic(46),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(155),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(161),
    to_slogic(156),
    to_slogic(165),
    to_slogic(157),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(143),
    to_slogic(135),
    to_slogic(121),
    to_slogic(100),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(134),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(135),
    to_slogic(126),
    to_slogic(134),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(134),
    to_slogic(130),
    to_slogic(126),
    to_slogic(134),
    to_slogic(130),
    to_slogic(133),
    to_slogic(128),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(124),
    to_slogic(116),
    to_slogic(124),
    to_slogic(121),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(128),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(119),
    to_slogic(118),
    to_slogic(117),
    to_slogic(116),
    to_slogic(110),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(128),
    to_slogic(142),
    to_slogic(137),
    to_slogic(146),
    to_slogic(152),
    to_slogic(155),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(158),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(156),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(143),
    to_slogic(144),
    to_slogic(136),
    to_slogic(144),
    to_slogic(172),
    to_slogic(196),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(222),
    to_slogic(213),
    to_slogic(183),
    to_slogic(125),
    to_slogic(109),
    to_slogic(101),
    to_slogic(116),
    to_slogic(107),
    to_slogic(116),
    to_slogic(117),
    to_slogic(126),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(99),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(42),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(100),
    to_slogic(89),
    to_slogic(82),
    to_slogic(92),
    to_slogic(94),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(121),
    to_slogic(117),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(124),
    to_slogic(128),
    to_slogic(134),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(118),
    to_slogic(121),
    to_slogic(121),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(128),
    to_slogic(126),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(119),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(146),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(183),
    to_slogic(207),
    to_slogic(213),
    to_slogic(222),
    to_slogic(223),
    to_slogic(222),
    to_slogic(213),
    to_slogic(197),
    to_slogic(158),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(124),
    to_slogic(133),
    to_slogic(126),
    to_slogic(94),
    to_slogic(49),
    to_slogic(44),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(155),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(151),
    to_slogic(143),
    to_slogic(135),
    to_slogic(121),
    to_slogic(99),
    to_slogic(89),
    to_slogic(81),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(117),
    to_slogic(116),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(126),
    to_slogic(121),
    to_slogic(128),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(121),
    to_slogic(117),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(116),
    to_slogic(121),
    to_slogic(121),
    to_slogic(117),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(128),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(117),
    to_slogic(126),
    to_slogic(124),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(103),
    to_slogic(109),
    to_slogic(119),
    to_slogic(128),
    to_slogic(133),
    to_slogic(137),
    to_slogic(146),
    to_slogic(143),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(136),
    to_slogic(144),
    to_slogic(165),
    to_slogic(197),
    to_slogic(213),
    to_slogic(222),
    to_slogic(223),
    to_slogic(223),
    to_slogic(222),
    to_slogic(213),
    to_slogic(191),
    to_slogic(136),
    to_slogic(94),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(117),
    to_slogic(92),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(97),
    to_slogic(82),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(121),
    to_slogic(117),
    to_slogic(124),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(117),
    to_slogic(130),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(128),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(124),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(121),
    to_slogic(124),
    to_slogic(126),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(116),
    to_slogic(121),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(124),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(126),
    to_slogic(128),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(119),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(150),
    to_slogic(152),
    to_slogic(155),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(184),
    to_slogic(205),
    to_slogic(213),
    to_slogic(222),
    to_slogic(223),
    to_slogic(223),
    to_slogic(222),
    to_slogic(205),
    to_slogic(172),
    to_slogic(107),
    to_slogic(109),
    to_slogic(107),
    to_slogic(109),
    to_slogic(117),
    to_slogic(116),
    to_slogic(107),
    to_slogic(128),
    to_slogic(118),
    to_slogic(133),
    to_slogic(126),
    to_slogic(92),
    to_slogic(56),
    to_slogic(44),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(161),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(165),
    to_slogic(156),
    to_slogic(157),
    to_slogic(157),
    to_slogic(161),
    to_slogic(157),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(116),
    to_slogic(99),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(116),
    to_slogic(117),
    to_slogic(126),
    to_slogic(118),
    to_slogic(124),
    to_slogic(126),
    to_slogic(121),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(121),
    to_slogic(124),
    to_slogic(121),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(121),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(124),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(117),
    to_slogic(134),
    to_slogic(128),
    to_slogic(128),
    to_slogic(124),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(130),
    to_slogic(128),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(110),
    to_slogic(109),
    to_slogic(109),
    to_slogic(118),
    to_slogic(119),
    to_slogic(119),
    to_slogic(134),
    to_slogic(137),
    to_slogic(137),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(155),
    to_slogic(152),
    to_slogic(157),
    to_slogic(155),
    to_slogic(152),
    to_slogic(156),
    to_slogic(157),
    to_slogic(144),
    to_slogic(157),
    to_slogic(152),
    to_slogic(150),
    to_slogic(156),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(136),
    to_slogic(143),
    to_slogic(143),
    to_slogic(165),
    to_slogic(191),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(223),
    to_slogic(222),
    to_slogic(213),
    to_slogic(197),
    to_slogic(136),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(117),
    to_slogic(118),
    to_slogic(133),
    to_slogic(126),
    to_slogic(89),
    to_slogic(63),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(156),
    to_slogic(151),
    to_slogic(151),
    to_slogic(156),
    to_slogic(151),
    to_slogic(156),
    to_slogic(161),
    to_slogic(157),
    to_slogic(156),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(151),
    to_slogic(151),
    to_slogic(130),
    to_slogic(109),
    to_slogic(100),
    to_slogic(82),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(121),
    to_slogic(116),
    to_slogic(121),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(128),
    to_slogic(124),
    to_slogic(134),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(130),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(134),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(141),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(143),
    to_slogic(141),
    to_slogic(139),
    to_slogic(125),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(121),
    to_slogic(126),
    to_slogic(119),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(109),
    to_slogic(119),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(110),
    to_slogic(109),
    to_slogic(128),
    to_slogic(128),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(143),
    to_slogic(144),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(155),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(156),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(184),
    to_slogic(205),
    to_slogic(213),
    to_slogic(222),
    to_slogic(223),
    to_slogic(223),
    to_slogic(222),
    to_slogic(205),
    to_slogic(176),
    to_slogic(107),
    to_slogic(102),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(107),
    to_slogic(94),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(156),
    to_slogic(151),
    to_slogic(156),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(143),
    to_slogic(135),
    to_slogic(117),
    to_slogic(100),
    to_slogic(92),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(116),
    to_slogic(126),
    to_slogic(117),
    to_slogic(126),
    to_slogic(124),
    to_slogic(121),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(134),
    to_slogic(128),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(133),
    to_slogic(134),
    to_slogic(141),
    to_slogic(144),
    to_slogic(141),
    to_slogic(144),
    to_slogic(149),
    to_slogic(165),
    to_slogic(167),
    to_slogic(170),
    to_slogic(176),
    to_slogic(170),
    to_slogic(182),
    to_slogic(176),
    to_slogic(185),
    to_slogic(177),
    to_slogic(170),
    to_slogic(156),
    to_slogic(132),
    to_slogic(128),
    to_slogic(117),
    to_slogic(116),
    to_slogic(116),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(119),
    to_slogic(117),
    to_slogic(109),
    to_slogic(119),
    to_slogic(109),
    to_slogic(118),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(126),
    to_slogic(134),
    to_slogic(137),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(155),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(156),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(156),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(137),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(144),
    to_slogic(157),
    to_slogic(191),
    to_slogic(213),
    to_slogic(213),
    to_slogic(223),
    to_slogic(222),
    to_slogic(222),
    to_slogic(222),
    to_slogic(197),
    to_slogic(143),
    to_slogic(116),
    to_slogic(107),
    to_slogic(107),
    to_slogic(117),
    to_slogic(117),
    to_slogic(118),
    to_slogic(92),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(151),
    to_slogic(156),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(156),
    to_slogic(143),
    to_slogic(135),
    to_slogic(121),
    to_slogic(97),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(97),
    to_slogic(99),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(94),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(124),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(128),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(128),
    to_slogic(124),
    to_slogic(128),
    to_slogic(135),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(134),
    to_slogic(141),
    to_slogic(151),
    to_slogic(142),
    to_slogic(149),
    to_slogic(155),
    to_slogic(144),
    to_slogic(143),
    to_slogic(157),
    to_slogic(165),
    to_slogic(167),
    to_slogic(162),
    to_slogic(176),
    to_slogic(170),
    to_slogic(182),
    to_slogic(177),
    to_slogic(170),
    to_slogic(185),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(185),
    to_slogic(189),
    to_slogic(176),
    to_slogic(158),
    to_slogic(141),
    to_slogic(118),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(126),
    to_slogic(128),
    to_slogic(133),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(117),
    to_slogic(115),
    to_slogic(109),
    to_slogic(118),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(133),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(137),
    to_slogic(144),
    to_slogic(152),
    to_slogic(139),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(150),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(156),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(152),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(144),
    to_slogic(136),
    to_slogic(144),
    to_slogic(144),
    to_slogic(172),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(223),
    to_slogic(223),
    to_slogic(222),
    to_slogic(222),
    to_slogic(184),
    to_slogic(124),
    to_slogic(109),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(92),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(46),
    to_slogic(40),
    to_slogic(44),
    to_slogic(46),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(161),
    to_slogic(156),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(135),
    to_slogic(143),
    to_slogic(151),
    to_slogic(157),
    to_slogic(161),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(165),
    to_slogic(157),
    to_slogic(161),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(121),
    to_slogic(100),
    to_slogic(81),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(124),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(128),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(127),
    to_slogic(141),
    to_slogic(144),
    to_slogic(143),
    to_slogic(157),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(149),
    to_slogic(172),
    to_slogic(170),
    to_slogic(172),
    to_slogic(165),
    to_slogic(170),
    to_slogic(176),
    to_slogic(185),
    to_slogic(176),
    to_slogic(176),
    to_slogic(182),
    to_slogic(171),
    to_slogic(170),
    to_slogic(176),
    to_slogic(182),
    to_slogic(189),
    to_slogic(176),
    to_slogic(189),
    to_slogic(189),
    to_slogic(176),
    to_slogic(156),
    to_slogic(125),
    to_slogic(117),
    to_slogic(116),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(119),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(124),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(109),
    to_slogic(110),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(117),
    to_slogic(124),
    to_slogic(133),
    to_slogic(139),
    to_slogic(137),
    to_slogic(152),
    to_slogic(144),
    to_slogic(146),
    to_slogic(137),
    to_slogic(152),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(156),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(143),
    to_slogic(137),
    to_slogic(151),
    to_slogic(183),
    to_slogic(205),
    to_slogic(213),
    to_slogic(223),
    to_slogic(223),
    to_slogic(223),
    to_slogic(223),
    to_slogic(205),
    to_slogic(165),
    to_slogic(118),
    to_slogic(117),
    to_slogic(116),
    to_slogic(96),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(157),
    to_slogic(165),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(151),
    to_slogic(143),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(143),
    to_slogic(151),
    to_slogic(156),
    to_slogic(165),
    to_slogic(161),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(161),
    to_slogic(152),
    to_slogic(143),
    to_slogic(135),
    to_slogic(109),
    to_slogic(97),
    to_slogic(81),
    to_slogic(89),
    to_slogic(89),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(115),
    to_slogic(109),
    to_slogic(117),
    to_slogic(116),
    to_slogic(118),
    to_slogic(116),
    to_slogic(124),
    to_slogic(121),
    to_slogic(117),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(121),
    to_slogic(124),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(128),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(124),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(124),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(151),
    to_slogic(141),
    to_slogic(142),
    to_slogic(151),
    to_slogic(149),
    to_slogic(141),
    to_slogic(141),
    to_slogic(144),
    to_slogic(149),
    to_slogic(155),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(165),
    to_slogic(172),
    to_slogic(176),
    to_slogic(176),
    to_slogic(185),
    to_slogic(176),
    to_slogic(170),
    to_slogic(170),
    to_slogic(170),
    to_slogic(182),
    to_slogic(176),
    to_slogic(176),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(158),
    to_slogic(128),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(128),
    to_slogic(119),
    to_slogic(124),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(117),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(102),
    to_slogic(110),
    to_slogic(117),
    to_slogic(119),
    to_slogic(133),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(139),
    to_slogic(151),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(143),
    to_slogic(139),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(130),
    to_slogic(144),
    to_slogic(143),
    to_slogic(158),
    to_slogic(197),
    to_slogic(213),
    to_slogic(222),
    to_slogic(223),
    to_slogic(223),
    to_slogic(223),
    to_slogic(222),
    to_slogic(205),
    to_slogic(144),
    to_slogic(117),
    to_slogic(94),
    to_slogic(63),
    to_slogic(40),
    to_slogic(46),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(156),
    to_slogic(143),
    to_slogic(135),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(157),
    to_slogic(161),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(156),
    to_slogic(143),
    to_slogic(135),
    to_slogic(121),
    to_slogic(92),
    to_slogic(81),
    to_slogic(82),
    to_slogic(81),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(116),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(130),
    to_slogic(121),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(128),
    to_slogic(130),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(128),
    to_slogic(134),
    to_slogic(134),
    to_slogic(141),
    to_slogic(134),
    to_slogic(127),
    to_slogic(125),
    to_slogic(141),
    to_slogic(144),
    to_slogic(141),
    to_slogic(144),
    to_slogic(144),
    to_slogic(141),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(149),
    to_slogic(143),
    to_slogic(151),
    to_slogic(158),
    to_slogic(162),
    to_slogic(156),
    to_slogic(167),
    to_slogic(158),
    to_slogic(176),
    to_slogic(182),
    to_slogic(170),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(171),
    to_slogic(176),
    to_slogic(183),
    to_slogic(176),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(200),
    to_slogic(193),
    to_slogic(177),
    to_slogic(144),
    to_slogic(117),
    to_slogic(116),
    to_slogic(116),
    to_slogic(119),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(124),
    to_slogic(128),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(118),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(126),
    to_slogic(134),
    to_slogic(144),
    to_slogic(137),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(144),
    to_slogic(151),
    to_slogic(151),
    to_slogic(143),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(139),
    to_slogic(143),
    to_slogic(139),
    to_slogic(136),
    to_slogic(135),
    to_slogic(144),
    to_slogic(136),
    to_slogic(144),
    to_slogic(136),
    to_slogic(143),
    to_slogic(144),
    to_slogic(130),
    to_slogic(144),
    to_slogic(184),
    to_slogic(205),
    to_slogic(213),
    to_slogic(223),
    to_slogic(223),
    to_slogic(223),
    to_slogic(223),
    to_slogic(222),
    to_slogic(183),
    to_slogic(116),
    to_slogic(63),
    to_slogic(44),
    to_slogic(42),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(121),
    to_slogic(109),
    to_slogic(135),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(161),
    to_slogic(157),
    to_slogic(156),
    to_slogic(151),
    to_slogic(135),
    to_slogic(109),
    to_slogic(97),
    to_slogic(81),
    to_slogic(75),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(115),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(121),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(121),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(125),
    to_slogic(128),
    to_slogic(119),
    to_slogic(125),
    to_slogic(133),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(151),
    to_slogic(149),
    to_slogic(151),
    to_slogic(149),
    to_slogic(151),
    to_slogic(158),
    to_slogic(149),
    to_slogic(158),
    to_slogic(172),
    to_slogic(165),
    to_slogic(167),
    to_slogic(165),
    to_slogic(171),
    to_slogic(167),
    to_slogic(176),
    to_slogic(176),
    to_slogic(170),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(193),
    to_slogic(189),
    to_slogic(193),
    to_slogic(193),
    to_slogic(196),
    to_slogic(193),
    to_slogic(193),
    to_slogic(158),
    to_slogic(120),
    to_slogic(109),
    to_slogic(118),
    to_slogic(119),
    to_slogic(124),
    to_slogic(119),
    to_slogic(126),
    to_slogic(117),
    to_slogic(124),
    to_slogic(119),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(116),
    to_slogic(109),
    to_slogic(117),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(118),
    to_slogic(124),
    to_slogic(128),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(151),
    to_slogic(139),
    to_slogic(152),
    to_slogic(152),
    to_slogic(150),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(151),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(135),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(135),
    to_slogic(156),
    to_slogic(191),
    to_slogic(213),
    to_slogic(222),
    to_slogic(223),
    to_slogic(223),
    to_slogic(223),
    to_slogic(223),
    to_slogic(205),
    to_slogic(94),
    to_slogic(42),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(115),
    to_slogic(97),
    to_slogic(121),
    to_slogic(130),
    to_slogic(144),
    to_slogic(151),
    to_slogic(156),
    to_slogic(172),
    to_slogic(161),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(156),
    to_slogic(156),
    to_slogic(143),
    to_slogic(135),
    to_slogic(121),
    to_slogic(97),
    to_slogic(81),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(96),
    to_slogic(102),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(124),
    to_slogic(121),
    to_slogic(126),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(124),
    to_slogic(128),
    to_slogic(121),
    to_slogic(128),
    to_slogic(124),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(139),
    to_slogic(125),
    to_slogic(125),
    to_slogic(127),
    to_slogic(117),
    to_slogic(119),
    to_slogic(127),
    to_slogic(125),
    to_slogic(139),
    to_slogic(132),
    to_slogic(134),
    to_slogic(125),
    to_slogic(134),
    to_slogic(141),
    to_slogic(134),
    to_slogic(139),
    to_slogic(143),
    to_slogic(155),
    to_slogic(149),
    to_slogic(151),
    to_slogic(158),
    to_slogic(167),
    to_slogic(158),
    to_slogic(165),
    to_slogic(167),
    to_slogic(165),
    to_slogic(170),
    to_slogic(170),
    to_slogic(182),
    to_slogic(176),
    to_slogic(176),
    to_slogic(189),
    to_slogic(182),
    to_slogic(193),
    to_slogic(183),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(193),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(185),
    to_slogic(141),
    to_slogic(119),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(115),
    to_slogic(115),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(116),
    to_slogic(119),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(152),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(136),
    to_slogic(139),
    to_slogic(136),
    to_slogic(143),
    to_slogic(144),
    to_slogic(136),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(135),
    to_slogic(144),
    to_slogic(172),
    to_slogic(197),
    to_slogic(213),
    to_slogic(223),
    to_slogic(223),
    to_slogic(223),
    to_slogic(222),
    to_slogic(196),
    to_slogic(70),
    to_slogic(40),
    to_slogic(40),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(97),
    to_slogic(97),
    to_slogic(109),
    to_slogic(135),
    to_slogic(151),
    to_slogic(156),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(151),
    to_slogic(143),
    to_slogic(135),
    to_slogic(115),
    to_slogic(97),
    to_slogic(81),
    to_slogic(75),
    to_slogic(81),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(115),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(124),
    to_slogic(121),
    to_slogic(126),
    to_slogic(117),
    to_slogic(121),
    to_slogic(124),
    to_slogic(126),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(121),
    to_slogic(124),
    to_slogic(130),
    to_slogic(162),
    to_slogic(124),
    to_slogic(128),
    to_slogic(128),
    to_slogic(125),
    to_slogic(128),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(120),
    to_slogic(128),
    to_slogic(120),
    to_slogic(134),
    to_slogic(132),
    to_slogic(134),
    to_slogic(134),
    to_slogic(125),
    to_slogic(139),
    to_slogic(141),
    to_slogic(133),
    to_slogic(139),
    to_slogic(151),
    to_slogic(144),
    to_slogic(151),
    to_slogic(158),
    to_slogic(158),
    to_slogic(158),
    to_slogic(157),
    to_slogic(167),
    to_slogic(158),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(189),
    to_slogic(189),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(189),
    to_slogic(193),
    to_slogic(189),
    to_slogic(193),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(200),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(153),
    to_slogic(119),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(124),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(126),
    to_slogic(134),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(146),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(191),
    to_slogic(207),
    to_slogic(223),
    to_slogic(223),
    to_slogic(223),
    to_slogic(213),
    to_slogic(136),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(97),
    to_slogic(81),
    to_slogic(89),
    to_slogic(115),
    to_slogic(135),
    to_slogic(144),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(161),
    to_slogic(151),
    to_slogic(143),
    to_slogic(135),
    to_slogic(115),
    to_slogic(89),
    to_slogic(75),
    to_slogic(76),
    to_slogic(82),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(96),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(116),
    to_slogic(117),
    to_slogic(116),
    to_slogic(115),
    to_slogic(117),
    to_slogic(126),
    to_slogic(117),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(121),
    to_slogic(124),
    to_slogic(121),
    to_slogic(158),
    to_slogic(135),
    to_slogic(92),
    to_slogic(117),
    to_slogic(119),
    to_slogic(119),
    to_slogic(118),
    to_slogic(117),
    to_slogic(128),
    to_slogic(119),
    to_slogic(128),
    to_slogic(119),
    to_slogic(128),
    to_slogic(139),
    to_slogic(125),
    to_slogic(133),
    to_slogic(133),
    to_slogic(125),
    to_slogic(134),
    to_slogic(132),
    to_slogic(139),
    to_slogic(139),
    to_slogic(141),
    to_slogic(144),
    to_slogic(141),
    to_slogic(149),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(165),
    to_slogic(170),
    to_slogic(167),
    to_slogic(171),
    to_slogic(170),
    to_slogic(182),
    to_slogic(189),
    to_slogic(176),
    to_slogic(189),
    to_slogic(189),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(182),
    to_slogic(182),
    to_slogic(196),
    to_slogic(193),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(193),
    to_slogic(176),
    to_slogic(132),
    to_slogic(107),
    to_slogic(102),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(116),
    to_slogic(109),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(118),
    to_slogic(109),
    to_slogic(110),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(118),
    to_slogic(124),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(143),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(143),
    to_slogic(135),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(157),
    to_slogic(205),
    to_slogic(222),
    to_slogic(222),
    to_slogic(213),
    to_slogic(156),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(151),
    to_slogic(130),
    to_slogic(121),
    to_slogic(89),
    to_slogic(76),
    to_slogic(89),
    to_slogic(109),
    to_slogic(135),
    to_slogic(143),
    to_slogic(156),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(156),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(115),
    to_slogic(89),
    to_slogic(81),
    to_slogic(76),
    to_slogic(75),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(102),
    to_slogic(99),
    to_slogic(96),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(116),
    to_slogic(115),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(117),
    to_slogic(121),
    to_slogic(124),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(151),
    to_slogic(116),
    to_slogic(109),
    to_slogic(119),
    to_slogic(117),
    to_slogic(128),
    to_slogic(117),
    to_slogic(119),
    to_slogic(127),
    to_slogic(118),
    to_slogic(119),
    to_slogic(119),
    to_slogic(125),
    to_slogic(128),
    to_slogic(134),
    to_slogic(125),
    to_slogic(125),
    to_slogic(125),
    to_slogic(134),
    to_slogic(134),
    to_slogic(137),
    to_slogic(133),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(149),
    to_slogic(149),
    to_slogic(165),
    to_slogic(167),
    to_slogic(170),
    to_slogic(182),
    to_slogic(170),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(193),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(193),
    to_slogic(158),
    to_slogic(107),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(110),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(110),
    to_slogic(124),
    to_slogic(133),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(137),
    to_slogic(137),
    to_slogic(144),
    to_slogic(137),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(183),
    to_slogic(213),
    to_slogic(205),
    to_slogic(158),
    to_slogic(70),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(33),
    to_slogic(33),
    to_slogic(173),
    to_slogic(172),
    to_slogic(165),
    to_slogic(161),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(100),
    to_slogic(76),
    to_slogic(75),
    to_slogic(89),
    to_slogic(121),
    to_slogic(135),
    to_slogic(143),
    to_slogic(151),
    to_slogic(161),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(157),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(116),
    to_slogic(89),
    to_slogic(76),
    to_slogic(76),
    to_slogic(82),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(96),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(94),
    to_slogic(102),
    to_slogic(94),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(116),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(116),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(143),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(127),
    to_slogic(130),
    to_slogic(137),
    to_slogic(125),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(125),
    to_slogic(127),
    to_slogic(141),
    to_slogic(132),
    to_slogic(134),
    to_slogic(144),
    to_slogic(151),
    to_slogic(155),
    to_slogic(158),
    to_slogic(167),
    to_slogic(167),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(182),
    to_slogic(177),
    to_slogic(182),
    to_slogic(182),
    to_slogic(185),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(193),
    to_slogic(196),
    to_slogic(200),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(193),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(196),
    to_slogic(165),
    to_slogic(109),
    to_slogic(96),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(110),
    to_slogic(92),
    to_slogic(102),
    to_slogic(109),
    to_slogic(124),
    to_slogic(134),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(146),
    to_slogic(152),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(133),
    to_slogic(139),
    to_slogic(137),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(152),
    to_slogic(157),
    to_slogic(165),
    to_slogic(191),
    to_slogic(143),
    to_slogic(64),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(63),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(173),
    to_slogic(172),
    to_slogic(161),
    to_slogic(152),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(89),
    to_slogic(76),
    to_slogic(76),
    to_slogic(99),
    to_slogic(109),
    to_slogic(130),
    to_slogic(143),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(115),
    to_slogic(89),
    to_slogic(76),
    to_slogic(70),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(96),
    to_slogic(92),
    to_slogic(101),
    to_slogic(102),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(94),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(115),
    to_slogic(116),
    to_slogic(124),
    to_slogic(116),
    to_slogic(121),
    to_slogic(124),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(121),
    to_slogic(124),
    to_slogic(116),
    to_slogic(144),
    to_slogic(133),
    to_slogic(109),
    to_slogic(117),
    to_slogic(116),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(119),
    to_slogic(119),
    to_slogic(128),
    to_slogic(127),
    to_slogic(118),
    to_slogic(133),
    to_slogic(127),
    to_slogic(128),
    to_slogic(125),
    to_slogic(139),
    to_slogic(125),
    to_slogic(146),
    to_slogic(133),
    to_slogic(134),
    to_slogic(134),
    to_slogic(132),
    to_slogic(139),
    to_slogic(139),
    to_slogic(151),
    to_slogic(144),
    to_slogic(149),
    to_slogic(157),
    to_slogic(158),
    to_slogic(167),
    to_slogic(167),
    to_slogic(171),
    to_slogic(167),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(193),
    to_slogic(189),
    to_slogic(196),
    to_slogic(193),
    to_slogic(189),
    to_slogic(196),
    to_slogic(196),
    to_slogic(193),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(193),
    to_slogic(176),
    to_slogic(109),
    to_slogic(88),
    to_slogic(94),
    to_slogic(94),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(119),
    to_slogic(139),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(128),
    to_slogic(133),
    to_slogic(134),
    to_slogic(126),
    to_slogic(134),
    to_slogic(139),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(121),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(68),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(96),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(99),
    to_slogic(81),
    to_slogic(81),
    to_slogic(81),
    to_slogic(92),
    to_slogic(116),
    to_slogic(130),
    to_slogic(151),
    to_slogic(151),
    to_slogic(165),
    to_slogic(169),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(121),
    to_slogic(89),
    to_slogic(76),
    to_slogic(76),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(96),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(115),
    to_slogic(116),
    to_slogic(117),
    to_slogic(116),
    to_slogic(124),
    to_slogic(116),
    to_slogic(121),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(121),
    to_slogic(121),
    to_slogic(124),
    to_slogic(130),
    to_slogic(165),
    to_slogic(116),
    to_slogic(115),
    to_slogic(116),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(118),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(125),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(137),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(141),
    to_slogic(149),
    to_slogic(144),
    to_slogic(155),
    to_slogic(149),
    to_slogic(166),
    to_slogic(158),
    to_slogic(165),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(185),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(200),
    to_slogic(193),
    to_slogic(196),
    to_slogic(193),
    to_slogic(189),
    to_slogic(196),
    to_slogic(196),
    to_slogic(189),
    to_slogic(191),
    to_slogic(196),
    to_slogic(197),
    to_slogic(208),
    to_slogic(192),
    to_slogic(170),
    to_slogic(149),
    to_slogic(96),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(103),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(118),
    to_slogic(117),
    to_slogic(139),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(139),
    to_slogic(134),
    to_slogic(128),
    to_slogic(119),
    to_slogic(116),
    to_slogic(128),
    to_slogic(128),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(135),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(126),
    to_slogic(70),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(83),
    to_slogic(146),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(81),
    to_slogic(82),
    to_slogic(82),
    to_slogic(81),
    to_slogic(99),
    to_slogic(116),
    to_slogic(130),
    to_slogic(143),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(89),
    to_slogic(76),
    to_slogic(75),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(103),
    to_slogic(96),
    to_slogic(99),
    to_slogic(102),
    to_slogic(92),
    to_slogic(96),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(117),
    to_slogic(116),
    to_slogic(115),
    to_slogic(109),
    to_slogic(116),
    to_slogic(124),
    to_slogic(116),
    to_slogic(121),
    to_slogic(117),
    to_slogic(124),
    to_slogic(121),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(135),
    to_slogic(144),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(119),
    to_slogic(118),
    to_slogic(133),
    to_slogic(125),
    to_slogic(125),
    to_slogic(128),
    to_slogic(137),
    to_slogic(132),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(144),
    to_slogic(151),
    to_slogic(143),
    to_slogic(151),
    to_slogic(158),
    to_slogic(158),
    to_slogic(172),
    to_slogic(171),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(182),
    to_slogic(196),
    to_slogic(196),
    to_slogic(189),
    to_slogic(193),
    to_slogic(196),
    to_slogic(189),
    to_slogic(191),
    to_slogic(196),
    to_slogic(205),
    to_slogic(208),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(220),
    to_slogic(165),
    to_slogic(82),
    to_slogic(92),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(110),
    to_slogic(126),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(128),
    to_slogic(121),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(124),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(143),
    to_slogic(139),
    to_slogic(144),
    to_slogic(143),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(143),
    to_slogic(82),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(83),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(68),
    to_slogic(133),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(116),
    to_slogic(99),
    to_slogic(81),
    to_slogic(89),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(121),
    to_slogic(135),
    to_slogic(151),
    to_slogic(151),
    to_slogic(161),
    to_slogic(165),
    to_slogic(169),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(92),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(99),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(96),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(135),
    to_slogic(121),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(133),
    to_slogic(125),
    to_slogic(128),
    to_slogic(128),
    to_slogic(127),
    to_slogic(134),
    to_slogic(134),
    to_slogic(133),
    to_slogic(139),
    to_slogic(125),
    to_slogic(139),
    to_slogic(132),
    to_slogic(151),
    to_slogic(139),
    to_slogic(151),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(171),
    to_slogic(176),
    to_slogic(176),
    to_slogic(189),
    to_slogic(189),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(182),
    to_slogic(191),
    to_slogic(189),
    to_slogic(193),
    to_slogic(189),
    to_slogic(196),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(177),
    to_slogic(191),
    to_slogic(208),
    to_slogic(208),
    to_slogic(208),
    to_slogic(220),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(220),
    to_slogic(125),
    to_slogic(82),
    to_slogic(89),
    to_slogic(100),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(103),
    to_slogic(102),
    to_slogic(109),
    to_slogic(117),
    to_slogic(134),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(156),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(130),
    to_slogic(116),
    to_slogic(100),
    to_slogic(99),
    to_slogic(102),
    to_slogic(117),
    to_slogic(126),
    to_slogic(139),
    to_slogic(146),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(102),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(68),
    to_slogic(81),
    to_slogic(56),
    to_slogic(40),
    to_slogic(75),
    to_slogic(120),
    to_slogic(150),
    to_slogic(162),
    to_slogic(157),
    to_slogic(156),
    to_slogic(143),
    to_slogic(121),
    to_slogic(109),
    to_slogic(81),
    to_slogic(82),
    to_slogic(89),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(116),
    to_slogic(130),
    to_slogic(144),
    to_slogic(156),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(115),
    to_slogic(89),
    to_slogic(81),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(94),
    to_slogic(102),
    to_slogic(100),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(116),
    to_slogic(115),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(126),
    to_slogic(117),
    to_slogic(121),
    to_slogic(121),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(119),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(117),
    to_slogic(128),
    to_slogic(119),
    to_slogic(117),
    to_slogic(128),
    to_slogic(119),
    to_slogic(124),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(128),
    to_slogic(133),
    to_slogic(134),
    to_slogic(133),
    to_slogic(134),
    to_slogic(139),
    to_slogic(146),
    to_slogic(134),
    to_slogic(137),
    to_slogic(149),
    to_slogic(155),
    to_slogic(158),
    to_slogic(167),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(185),
    to_slogic(185),
    to_slogic(189),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(182),
    to_slogic(176),
    to_slogic(185),
    to_slogic(191),
    to_slogic(208),
    to_slogic(208),
    to_slogic(214),
    to_slogic(213),
    to_slogic(208),
    to_slogic(214),
    to_slogic(214),
    to_slogic(208),
    to_slogic(213),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(226),
    to_slogic(177),
    to_slogic(96),
    to_slogic(82),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(96),
    to_slogic(102),
    to_slogic(96),
    to_slogic(92),
    to_slogic(102),
    to_slogic(110),
    to_slogic(126),
    to_slogic(133),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(134),
    to_slogic(117),
    to_slogic(99),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(118),
    to_slogic(133),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(121),
    to_slogic(63),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(68),
    to_slogic(83),
    to_slogic(63),
    to_slogic(49),
    to_slogic(69),
    to_slogic(109),
    to_slogic(151),
    to_slogic(150),
    to_slogic(165),
    to_slogic(156),
    to_slogic(143),
    to_slogic(135),
    to_slogic(109),
    to_slogic(92),
    to_slogic(81),
    to_slogic(89),
    to_slogic(82),
    to_slogic(89),
    to_slogic(82),
    to_slogic(99),
    to_slogic(116),
    to_slogic(135),
    to_slogic(143),
    to_slogic(151),
    to_slogic(161),
    to_slogic(165),
    to_slogic(169),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(109),
    to_slogic(92),
    to_slogic(76),
    to_slogic(76),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(100),
    to_slogic(102),
    to_slogic(96),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(116),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(121),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(130),
    to_slogic(121),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(119),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(117),
    to_slogic(119),
    to_slogic(118),
    to_slogic(119),
    to_slogic(118),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(125),
    to_slogic(133),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(137),
    to_slogic(134),
    to_slogic(133),
    to_slogic(139),
    to_slogic(139),
    to_slogic(130),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(155),
    to_slogic(167),
    to_slogic(167),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(193),
    to_slogic(182),
    to_slogic(189),
    to_slogic(182),
    to_slogic(176),
    to_slogic(170),
    to_slogic(177),
    to_slogic(192),
    to_slogic(205),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(208),
    to_slogic(208),
    to_slogic(208),
    to_slogic(208),
    to_slogic(213),
    to_slogic(208),
    to_slogic(205),
    to_slogic(208),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(165),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(99),
    to_slogic(87),
    to_slogic(102),
    to_slogic(109),
    to_slogic(117),
    to_slogic(134),
    to_slogic(144),
    to_slogic(144),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(146),
    to_slogic(144),
    to_slogic(139),
    to_slogic(117),
    to_slogic(92),
    to_slogic(70),
    to_slogic(63),
    to_slogic(82),
    to_slogic(109),
    to_slogic(128),
    to_slogic(133),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(126),
    to_slogic(69),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(36),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(75),
    to_slogic(69),
    to_slogic(63),
    to_slogic(75),
    to_slogic(109),
    to_slogic(139),
    to_slogic(152),
    to_slogic(143),
    to_slogic(155),
    to_slogic(143),
    to_slogic(143),
    to_slogic(115),
    to_slogic(100),
    to_slogic(81),
    to_slogic(89),
    to_slogic(82),
    to_slogic(92),
    to_slogic(89),
    to_slogic(82),
    to_slogic(92),
    to_slogic(116),
    to_slogic(135),
    to_slogic(143),
    to_slogic(157),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(97),
    to_slogic(82),
    to_slogic(75),
    to_slogic(81),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(115),
    to_slogic(116),
    to_slogic(115),
    to_slogic(116),
    to_slogic(117),
    to_slogic(121),
    to_slogic(121),
    to_slogic(117),
    to_slogic(124),
    to_slogic(126),
    to_slogic(124),
    to_slogic(121),
    to_slogic(130),
    to_slogic(116),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(119),
    to_slogic(128),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(118),
    to_slogic(133),
    to_slogic(125),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(137),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(141),
    to_slogic(150),
    to_slogic(155),
    to_slogic(162),
    to_slogic(165),
    to_slogic(176),
    to_slogic(182),
    to_slogic(171),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(167),
    to_slogic(162),
    to_slogic(177),
    to_slogic(197),
    to_slogic(208),
    to_slogic(214),
    to_slogic(214),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(214),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(213),
    to_slogic(214),
    to_slogic(205),
    to_slogic(213),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(214),
    to_slogic(143),
    to_slogic(75),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(96),
    to_slogic(102),
    to_slogic(96),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(109),
    to_slogic(118),
    to_slogic(133),
    to_slogic(144),
    to_slogic(146),
    to_slogic(157),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(139),
    to_slogic(117),
    to_slogic(99),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(92),
    to_slogic(118),
    to_slogic(128),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(157),
    to_slogic(144),
    to_slogic(99),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(33),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(68),
    to_slogic(71),
    to_slogic(63),
    to_slogic(81),
    to_slogic(63),
    to_slogic(81),
    to_slogic(109),
    to_slogic(139),
    to_slogic(151),
    to_slogic(143),
    to_slogic(152),
    to_slogic(152),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(82),
    to_slogic(89),
    to_slogic(82),
    to_slogic(82),
    to_slogic(89),
    to_slogic(89),
    to_slogic(89),
    to_slogic(99),
    to_slogic(116),
    to_slogic(135),
    to_slogic(144),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(115),
    to_slogic(92),
    to_slogic(81),
    to_slogic(76),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(96),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(96),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(115),
    to_slogic(117),
    to_slogic(117),
    to_slogic(116),
    to_slogic(117),
    to_slogic(121),
    to_slogic(124),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(126),
    to_slogic(126),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(128),
    to_slogic(133),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(133),
    to_slogic(137),
    to_slogic(134),
    to_slogic(137),
    to_slogic(149),
    to_slogic(139),
    to_slogic(146),
    to_slogic(143),
    to_slogic(151),
    to_slogic(141),
    to_slogic(149),
    to_slogic(149),
    to_slogic(165),
    to_slogic(156),
    to_slogic(171),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(166),
    to_slogic(162),
    to_slogic(165),
    to_slogic(191),
    to_slogic(205),
    to_slogic(214),
    to_slogic(214),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(205),
    to_slogic(214),
    to_slogic(208),
    to_slogic(226),
    to_slogic(220),
    to_slogic(213),
    to_slogic(114),
    to_slogic(75),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(96),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(109),
    to_slogic(117),
    to_slogic(134),
    to_slogic(139),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(139),
    to_slogic(119),
    to_slogic(102),
    to_slogic(63),
    to_slogic(44),
    to_slogic(56),
    to_slogic(81),
    to_slogic(102),
    to_slogic(117),
    to_slogic(134),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(115),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(68),
    to_slogic(71),
    to_slogic(81),
    to_slogic(81),
    to_slogic(109),
    to_slogic(132),
    to_slogic(151),
    to_slogic(155),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(97),
    to_slogic(89),
    to_slogic(82),
    to_slogic(92),
    to_slogic(89),
    to_slogic(89),
    to_slogic(81),
    to_slogic(82),
    to_slogic(94),
    to_slogic(116),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(135),
    to_slogic(130),
    to_slogic(115),
    to_slogic(89),
    to_slogic(81),
    to_slogic(76),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(96),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(121),
    to_slogic(115),
    to_slogic(116),
    to_slogic(124),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(121),
    to_slogic(117),
    to_slogic(130),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(115),
    to_slogic(110),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(101),
    to_slogic(119),
    to_slogic(128),
    to_slogic(118),
    to_slogic(128),
    to_slogic(120),
    to_slogic(128),
    to_slogic(134),
    to_slogic(137),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(137),
    to_slogic(137),
    to_slogic(146),
    to_slogic(143),
    to_slogic(146),
    to_slogic(143),
    to_slogic(146),
    to_slogic(152),
    to_slogic(151),
    to_slogic(155),
    to_slogic(165),
    to_slogic(176),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(158),
    to_slogic(162),
    to_slogic(185),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(197),
    to_slogic(205),
    to_slogic(208),
    to_slogic(208),
    to_slogic(220),
    to_slogic(214),
    to_slogic(220),
    to_slogic(226),
    to_slogic(226),
    to_slogic(220),
    to_slogic(191),
    to_slogic(91),
    to_slogic(75),
    to_slogic(81),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(87),
    to_slogic(99),
    to_slogic(110),
    to_slogic(117),
    to_slogic(134),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(149),
    to_slogic(146),
    to_slogic(144),
    to_slogic(128),
    to_slogic(102),
    to_slogic(76),
    to_slogic(44),
    to_slogic(44),
    to_slogic(62),
    to_slogic(92),
    to_slogic(109),
    to_slogic(128),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(152),
    to_slogic(130),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(68),
    to_slogic(71),
    to_slogic(75),
    to_slogic(81),
    to_slogic(101),
    to_slogic(125),
    to_slogic(144),
    to_slogic(143),
    to_slogic(155),
    to_slogic(143),
    to_slogic(139),
    to_slogic(155),
    to_slogic(121),
    to_slogic(100),
    to_slogic(89),
    to_slogic(82),
    to_slogic(92),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(81),
    to_slogic(99),
    to_slogic(109),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(92),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(83),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(115),
    to_slogic(117),
    to_slogic(116),
    to_slogic(116),
    to_slogic(124),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(116),
    to_slogic(116),
    to_slogic(109),
    to_slogic(100),
    to_slogic(117),
    to_slogic(118),
    to_slogic(109),
    to_slogic(109),
    to_slogic(110),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(119),
    to_slogic(109),
    to_slogic(101),
    to_slogic(119),
    to_slogic(117),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(137),
    to_slogic(137),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(151),
    to_slogic(146),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(151),
    to_slogic(162),
    to_slogic(162),
    to_slogic(167),
    to_slogic(176),
    to_slogic(172),
    to_slogic(156),
    to_slogic(151),
    to_slogic(165),
    to_slogic(197),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(196),
    to_slogic(204),
    to_slogic(197),
    to_slogic(214),
    to_slogic(211),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(214),
    to_slogic(220),
    to_slogic(205),
    to_slogic(220),
    to_slogic(208),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(220),
    to_slogic(165),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(109),
    to_slogic(124),
    to_slogic(134),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(139),
    to_slogic(128),
    to_slogic(102),
    to_slogic(62),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(82),
    to_slogic(102),
    to_slogic(117),
    to_slogic(134),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(152),
    to_slogic(144),
    to_slogic(92),
    to_slogic(44),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(46),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(65),
    to_slogic(75),
    to_slogic(81),
    to_slogic(110),
    to_slogic(132),
    to_slogic(144),
    to_slogic(151),
    to_slogic(149),
    to_slogic(152),
    to_slogic(137),
    to_slogic(150),
    to_slogic(162),
    to_slogic(100),
    to_slogic(92),
    to_slogic(82),
    to_slogic(89),
    to_slogic(82),
    to_slogic(92),
    to_slogic(89),
    to_slogic(89),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(115),
    to_slogic(135),
    to_slogic(143),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(152),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(94),
    to_slogic(76),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(96),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(117),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(126),
    to_slogic(128),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(116),
    to_slogic(107),
    to_slogic(117),
    to_slogic(119),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(125),
    to_slogic(128),
    to_slogic(125),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(137),
    to_slogic(146),
    to_slogic(139),
    to_slogic(146),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(146),
    to_slogic(141),
    to_slogic(149),
    to_slogic(155),
    to_slogic(165),
    to_slogic(171),
    to_slogic(162),
    to_slogic(139),
    to_slogic(149),
    to_slogic(177),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(211),
    to_slogic(204),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(197),
    to_slogic(204),
    to_slogic(208),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(208),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(208),
    to_slogic(153),
    to_slogic(102),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(81),
    to_slogic(89),
    to_slogic(82),
    to_slogic(92),
    to_slogic(109),
    to_slogic(124),
    to_slogic(130),
    to_slogic(139),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(124),
    to_slogic(100),
    to_slogic(70),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(75),
    to_slogic(96),
    to_slogic(109),
    to_slogic(130),
    to_slogic(133),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(116),
    to_slogic(56),
    to_slogic(40),
    to_slogic(36),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(81),
    to_slogic(102),
    to_slogic(125),
    to_slogic(141),
    to_slogic(151),
    to_slogic(149),
    to_slogic(139),
    to_slogic(139),
    to_slogic(150),
    to_slogic(162),
    to_slogic(158),
    to_slogic(92),
    to_slogic(81),
    to_slogic(89),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(81),
    to_slogic(100),
    to_slogic(109),
    to_slogic(130),
    to_slogic(144),
    to_slogic(151),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(130),
    to_slogic(115),
    to_slogic(92),
    to_slogic(75),
    to_slogic(70),
    to_slogic(76),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(102),
    to_slogic(94),
    to_slogic(102),
    to_slogic(102),
    to_slogic(99),
    to_slogic(96),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(121),
    to_slogic(117),
    to_slogic(116),
    to_slogic(116),
    to_slogic(118),
    to_slogic(116),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(133),
    to_slogic(116),
    to_slogic(115),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(119),
    to_slogic(117),
    to_slogic(119),
    to_slogic(128),
    to_slogic(124),
    to_slogic(128),
    to_slogic(134),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(137),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(137),
    to_slogic(134),
    to_slogic(146),
    to_slogic(139),
    to_slogic(152),
    to_slogic(149),
    to_slogic(155),
    to_slogic(166),
    to_slogic(155),
    to_slogic(132),
    to_slogic(155),
    to_slogic(189),
    to_slogic(191),
    to_slogic(200),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(211),
    to_slogic(197),
    to_slogic(196),
    to_slogic(205),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(208),
    to_slogic(208),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(226),
    to_slogic(196),
    to_slogic(133),
    to_slogic(75),
    to_slogic(70),
    to_slogic(75),
    to_slogic(89),
    to_slogic(82),
    to_slogic(92),
    to_slogic(102),
    to_slogic(116),
    to_slogic(134),
    to_slogic(144),
    to_slogic(144),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(139),
    to_slogic(126),
    to_slogic(94),
    to_slogic(76),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(76),
    to_slogic(99),
    to_slogic(117),
    to_slogic(130),
    to_slogic(139),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(151),
    to_slogic(130),
    to_slogic(76),
    to_slogic(44),
    to_slogic(40),
    to_slogic(36),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(96),
    to_slogic(125),
    to_slogic(143),
    to_slogic(151),
    to_slogic(144),
    to_slogic(151),
    to_slogic(143),
    to_slogic(149),
    to_slogic(158),
    to_slogic(166),
    to_slogic(162),
    to_slogic(92),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(109),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(144),
    to_slogic(121),
    to_slogic(116),
    to_slogic(99),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(89),
    to_slogic(92),
    to_slogic(99),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(92),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(115),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(124),
    to_slogic(116),
    to_slogic(126),
    to_slogic(135),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(110),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(125),
    to_slogic(133),
    to_slogic(134),
    to_slogic(128),
    to_slogic(125),
    to_slogic(133),
    to_slogic(139),
    to_slogic(146),
    to_slogic(133),
    to_slogic(137),
    to_slogic(146),
    to_slogic(139),
    to_slogic(146),
    to_slogic(133),
    to_slogic(139),
    to_slogic(125),
    to_slogic(133),
    to_slogic(139),
    to_slogic(137),
    to_slogic(141),
    to_slogic(143),
    to_slogic(155),
    to_slogic(151),
    to_slogic(141),
    to_slogic(170),
    to_slogic(196),
    to_slogic(191),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(208),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(205),
    to_slogic(208),
    to_slogic(208),
    to_slogic(208),
    to_slogic(208),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(208),
    to_slogic(149),
    to_slogic(75),
    to_slogic(70),
    to_slogic(76),
    to_slogic(75),
    to_slogic(92),
    to_slogic(100),
    to_slogic(124),
    to_slogic(134),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(149),
    to_slogic(144),
    to_slogic(124),
    to_slogic(100),
    to_slogic(76),
    to_slogic(44),
    to_slogic(49),
    to_slogic(33),
    to_slogic(44),
    to_slogic(56),
    to_slogic(81),
    to_slogic(102),
    to_slogic(124),
    to_slogic(133),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(99),
    to_slogic(44),
    to_slogic(33),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(81),
    to_slogic(120),
    to_slogic(141),
    to_slogic(141),
    to_slogic(143),
    to_slogic(151),
    to_slogic(143),
    to_slogic(144),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(82),
    to_slogic(102),
    to_slogic(109),
    to_slogic(130),
    to_slogic(144),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(115),
    to_slogic(92),
    to_slogic(81),
    to_slogic(76),
    to_slogic(75),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(94),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(116),
    to_slogic(117),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(143),
    to_slogic(116),
    to_slogic(115),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(146),
    to_slogic(139),
    to_slogic(146),
    to_slogic(134),
    to_slogic(146),
    to_slogic(134),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(146),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(144),
    to_slogic(182),
    to_slogic(189),
    to_slogic(200),
    to_slogic(196),
    to_slogic(196),
    to_slogic(193),
    to_slogic(196),
    to_slogic(189),
    to_slogic(196),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(200),
    to_slogic(196),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(205),
    to_slogic(205),
    to_slogic(213),
    to_slogic(208),
    to_slogic(213),
    to_slogic(205),
    to_slogic(214),
    to_slogic(214),
    to_slogic(205),
    to_slogic(220),
    to_slogic(226),
    to_slogic(208),
    to_slogic(109),
    to_slogic(56),
    to_slogic(70),
    to_slogic(70),
    to_slogic(92),
    to_slogic(102),
    to_slogic(117),
    to_slogic(130),
    to_slogic(139),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(144),
    to_slogic(139),
    to_slogic(117),
    to_slogic(102),
    to_slogic(76),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(62),
    to_slogic(89),
    to_slogic(109),
    to_slogic(126),
    to_slogic(139),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(117),
    to_slogic(56),
    to_slogic(44),
    to_slogic(40),
    to_slogic(46),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(56),
    to_slogic(81),
    to_slogic(120),
    to_slogic(141),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(143),
    to_slogic(156),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(82),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(116),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(143),
    to_slogic(130),
    to_slogic(116),
    to_slogic(92),
    to_slogic(82),
    to_slogic(77),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(116),
    to_slogic(115),
    to_slogic(150),
    to_slogic(144),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(118),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(152),
    to_slogic(139),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(146),
    to_slogic(141),
    to_slogic(139),
    to_slogic(146),
    to_slogic(133),
    to_slogic(134),
    to_slogic(133),
    to_slogic(127),
    to_slogic(137),
    to_slogic(125),
    to_slogic(128),
    to_slogic(141),
    to_slogic(165),
    to_slogic(176),
    to_slogic(182),
    to_slogic(189),
    to_slogic(196),
    to_slogic(200),
    to_slogic(196),
    to_slogic(189),
    to_slogic(193),
    to_slogic(191),
    to_slogic(185),
    to_slogic(196),
    to_slogic(191),
    to_slogic(193),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(211),
    to_slogic(204),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(213),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(208),
    to_slogic(208),
    to_slogic(213),
    to_slogic(214),
    to_slogic(220),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(193),
    to_slogic(82),
    to_slogic(62),
    to_slogic(76),
    to_slogic(81),
    to_slogic(94),
    to_slogic(117),
    to_slogic(130),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(149),
    to_slogic(157),
    to_slogic(152),
    to_slogic(146),
    to_slogic(144),
    to_slogic(124),
    to_slogic(109),
    to_slogic(75),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(33),
    to_slogic(44),
    to_slogic(56),
    to_slogic(76),
    to_slogic(97),
    to_slogic(116),
    to_slogic(130),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(130),
    to_slogic(75),
    to_slogic(44),
    to_slogic(40),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(68),
    to_slogic(110),
    to_slogic(141),
    to_slogic(144),
    to_slogic(151),
    to_slogic(139),
    to_slogic(139),
    to_slogic(141),
    to_slogic(156),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(82),
    to_slogic(99),
    to_slogic(116),
    to_slogic(130),
    to_slogic(143),
    to_slogic(152),
    to_slogic(152),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(144),
    to_slogic(126),
    to_slogic(115),
    to_slogic(92),
    to_slogic(82),
    to_slogic(75),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(96),
    to_slogic(99),
    to_slogic(102),
    to_slogic(96),
    to_slogic(100),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(117),
    to_slogic(116),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(117),
    to_slogic(178),
    to_slogic(135),
    to_slogic(99),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(119),
    to_slogic(133),
    to_slogic(134),
    to_slogic(133),
    to_slogic(139),
    to_slogic(146),
    to_slogic(137),
    to_slogic(128),
    to_slogic(137),
    to_slogic(137),
    to_slogic(139),
    to_slogic(146),
    to_slogic(139),
    to_slogic(133),
    to_slogic(133),
    to_slogic(125),
    to_slogic(128),
    to_slogic(124),
    to_slogic(128),
    to_slogic(127),
    to_slogic(144),
    to_slogic(171),
    to_slogic(189),
    to_slogic(182),
    to_slogic(182),
    to_slogic(193),
    to_slogic(195),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(191),
    to_slogic(189),
    to_slogic(196),
    to_slogic(185),
    to_slogic(185),
    to_slogic(185),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(208),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(133),
    to_slogic(75),
    to_slogic(63),
    to_slogic(81),
    to_slogic(92),
    to_slogic(115),
    to_slogic(130),
    to_slogic(139),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(146),
    to_slogic(139),
    to_slogic(126),
    to_slogic(102),
    to_slogic(75),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(33),
    to_slogic(33),
    to_slogic(56),
    to_slogic(81),
    to_slogic(100),
    to_slogic(121),
    to_slogic(130),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(135),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(100),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(65),
    to_slogic(101),
    to_slogic(133),
    to_slogic(149),
    to_slogic(152),
    to_slogic(141),
    to_slogic(132),
    to_slogic(139),
    to_slogic(149),
    to_slogic(158),
    to_slogic(162),
    to_slogic(162),
    to_slogic(158),
    to_slogic(166),
    to_slogic(162),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(109),
    to_slogic(130),
    to_slogic(144),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(152),
    to_slogic(144),
    to_slogic(130),
    to_slogic(116),
    to_slogic(92),
    to_slogic(82),
    to_slogic(77),
    to_slogic(82),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(115),
    to_slogic(115),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(144),
    to_slogic(183),
    to_slogic(130),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(134),
    to_slogic(146),
    to_slogic(133),
    to_slogic(125),
    to_slogic(133),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(133),
    to_slogic(133),
    to_slogic(125),
    to_slogic(128),
    to_slogic(119),
    to_slogic(110),
    to_slogic(120),
    to_slogic(158),
    to_slogic(172),
    to_slogic(182),
    to_slogic(189),
    to_slogic(200),
    to_slogic(193),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(185),
    to_slogic(182),
    to_slogic(191),
    to_slogic(196),
    to_slogic(197),
    to_slogic(200),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(200),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(220),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(226),
    to_slogic(226),
    to_slogic(197),
    to_slogic(114),
    to_slogic(62),
    to_slogic(76),
    to_slogic(89),
    to_slogic(109),
    to_slogic(126),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(144),
    to_slogic(139),
    to_slogic(124),
    to_slogic(102),
    to_slogic(82),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(33),
    to_slogic(44),
    to_slogic(56),
    to_slogic(81),
    to_slogic(100),
    to_slogic(116),
    to_slogic(137),
    to_slogic(155),
    to_slogic(158),
    to_slogic(158),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(121),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(87),
    to_slogic(126),
    to_slogic(151),
    to_slogic(151),
    to_slogic(141),
    to_slogic(132),
    to_slogic(139),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(82),
    to_slogic(92),
    to_slogic(109),
    to_slogic(130),
    to_slogic(144),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(152),
    to_slogic(143),
    to_slogic(130),
    to_slogic(118),
    to_slogic(92),
    to_slogic(75),
    to_slogic(76),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(96),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(117),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(183),
    to_slogic(172),
    to_slogic(115),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(118),
    to_slogic(119),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(134),
    to_slogic(139),
    to_slogic(137),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(139),
    to_slogic(133),
    to_slogic(134),
    to_slogic(146),
    to_slogic(139),
    to_slogic(133),
    to_slogic(120),
    to_slogic(128),
    to_slogic(119),
    to_slogic(101),
    to_slogic(134),
    to_slogic(165),
    to_slogic(182),
    to_slogic(182),
    to_slogic(187),
    to_slogic(185),
    to_slogic(193),
    to_slogic(185),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(185),
    to_slogic(176),
    to_slogic(177),
    to_slogic(200),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(195),
    to_slogic(200),
    to_slogic(197),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(214),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(226),
    to_slogic(226),
    to_slogic(191),
    to_slogic(69),
    to_slogic(63),
    to_slogic(82),
    to_slogic(116),
    to_slogic(134),
    to_slogic(139),
    to_slogic(144),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(146),
    to_slogic(139),
    to_slogic(126),
    to_slogic(102),
    to_slogic(75),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(40),
    to_slogic(44),
    to_slogic(33),
    to_slogic(33),
    to_slogic(56),
    to_slogic(91),
    to_slogic(149),
    to_slogic(191),
    to_slogic(208),
    to_slogic(220),
    to_slogic(208),
    to_slogic(185),
    to_slogic(179),
    to_slogic(191),
    to_slogic(166),
    to_slogic(133),
    to_slogic(75),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(75),
    to_slogic(120),
    to_slogic(151),
    to_slogic(151),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(149),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(158),
    to_slogic(162),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(82),
    to_slogic(89),
    to_slogic(82),
    to_slogic(89),
    to_slogic(81),
    to_slogic(89),
    to_slogic(92),
    to_slogic(109),
    to_slogic(130),
    to_slogic(143),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(151),
    to_slogic(144),
    to_slogic(130),
    to_slogic(117),
    to_slogic(92),
    to_slogic(82),
    to_slogic(76),
    to_slogic(82),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(102),
    to_slogic(96),
    to_slogic(100),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(102),
    to_slogic(128),
    to_slogic(205),
    to_slogic(165),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(117),
    to_slogic(117),
    to_slogic(126),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(137),
    to_slogic(133),
    to_slogic(133),
    to_slogic(134),
    to_slogic(137),
    to_slogic(137),
    to_slogic(119),
    to_slogic(117),
    to_slogic(128),
    to_slogic(119),
    to_slogic(109),
    to_slogic(151),
    to_slogic(162),
    to_slogic(166),
    to_slogic(193),
    to_slogic(189),
    to_slogic(182),
    to_slogic(183),
    to_slogic(176),
    to_slogic(182),
    to_slogic(191),
    to_slogic(191),
    to_slogic(182),
    to_slogic(167),
    to_slogic(172),
    to_slogic(189),
    to_slogic(193),
    to_slogic(191),
    to_slogic(200),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(197),
    to_slogic(205),
    to_slogic(197),
    to_slogic(196),
    to_slogic(197),
    to_slogic(197),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(220),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(208),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(226),
    to_slogic(220),
    to_slogic(96),
    to_slogic(63),
    to_slogic(89),
    to_slogic(109),
    to_slogic(126),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(139),
    to_slogic(119),
    to_slogic(109),
    to_slogic(75),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(40),
    to_slogic(81),
    to_slogic(177),
    to_slogic(214),
    to_slogic(220),
    to_slogic(207),
    to_slogic(196),
    to_slogic(196),
    to_slogic(208),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(133),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(75),
    to_slogic(110),
    to_slogic(141),
    to_slogic(149),
    to_slogic(143),
    to_slogic(141),
    to_slogic(139),
    to_slogic(144),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(155),
    to_slogic(162),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(82),
    to_slogic(89),
    to_slogic(109),
    to_slogic(121),
    to_slogic(144),
    to_slogic(152),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(152),
    to_slogic(143),
    to_slogic(130),
    to_slogic(116),
    to_slogic(92),
    to_slogic(76),
    to_slogic(69),
    to_slogic(81),
    to_slogic(82),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(96),
    to_slogic(92),
    to_slogic(99),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(173),
    to_slogic(203),
    to_slogic(143),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(118),
    to_slogic(109),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(133),
    to_slogic(137),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(137),
    to_slogic(133),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(110),
    to_slogic(127),
    to_slogic(149),
    to_slogic(167),
    to_slogic(176),
    to_slogic(176),
    to_slogic(193),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(167),
    to_slogic(182),
    to_slogic(189),
    to_slogic(182),
    to_slogic(179),
    to_slogic(185),
    to_slogic(195),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(200),
    to_slogic(191),
    to_slogic(200),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(200),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(204),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(196),
    to_slogic(205),
    to_slogic(208),
    to_slogic(205),
    to_slogic(214),
    to_slogic(205),
    to_slogic(208),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(226),
    to_slogic(226),
    to_slogic(153),
    to_slogic(63),
    to_slogic(81),
    to_slogic(102),
    to_slogic(126),
    to_slogic(139),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(139),
    to_slogic(126),
    to_slogic(109),
    to_slogic(75),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(49),
    to_slogic(102),
    to_slogic(191),
    to_slogic(220),
    to_slogic(213),
    to_slogic(196),
    to_slogic(196),
    to_slogic(208),
    to_slogic(208),
    to_slogic(220),
    to_slogic(226),
    to_slogic(226),
    to_slogic(220),
    to_slogic(177),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(40),
    to_slogic(56),
    to_slogic(89),
    to_slogic(141),
    to_slogic(144),
    to_slogic(151),
    to_slogic(141),
    to_slogic(141),
    to_slogic(144),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(92),
    to_slogic(92),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(82),
    to_slogic(82),
    to_slogic(89),
    to_slogic(109),
    to_slogic(130),
    to_slogic(139),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(89),
    to_slogic(77),
    to_slogic(70),
    to_slogic(76),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(94),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(102),
    to_slogic(118),
    to_slogic(198),
    to_slogic(184),
    to_slogic(152),
    to_slogic(115),
    to_slogic(99),
    to_slogic(102),
    to_slogic(102),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(115),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(119),
    to_slogic(133),
    to_slogic(133),
    to_slogic(137),
    to_slogic(130),
    to_slogic(128),
    to_slogic(128),
    to_slogic(107),
    to_slogic(101),
    to_slogic(133),
    to_slogic(158),
    to_slogic(172),
    to_slogic(172),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(185),
    to_slogic(167),
    to_slogic(158),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(182),
    to_slogic(185),
    to_slogic(185),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(200),
    to_slogic(196),
    to_slogic(191),
    to_slogic(200),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(193),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(214),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(213),
    to_slogic(220),
    to_slogic(226),
    to_slogic(226),
    to_slogic(197),
    to_slogic(96),
    to_slogic(69),
    to_slogic(100),
    to_slogic(121),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(139),
    to_slogic(121),
    to_slogic(100),
    to_slogic(75),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(56),
    to_slogic(127),
    to_slogic(196),
    to_slogic(220),
    to_slogic(196),
    to_slogic(176),
    to_slogic(196),
    to_slogic(214),
    to_slogic(220),
    to_slogic(226),
    to_slogic(220),
    to_slogic(226),
    to_slogic(226),
    to_slogic(226),
    to_slogic(226),
    to_slogic(96),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(81),
    to_slogic(125),
    to_slogic(151),
    to_slogic(151),
    to_slogic(144),
    to_slogic(139),
    to_slogic(141),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(150),
    to_slogic(162),
    to_slogic(155),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(89),
    to_slogic(92),
    to_slogic(109),
    to_slogic(130),
    to_slogic(135),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(143),
    to_slogic(130),
    to_slogic(115),
    to_slogic(89),
    to_slogic(70),
    to_slogic(70),
    to_slogic(76),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(102),
    to_slogic(99),
    to_slogic(99),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(128),
    to_slogic(205),
    to_slogic(176),
    to_slogic(143),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(118),
    to_slogic(116),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(126),
    to_slogic(124),
    to_slogic(118),
    to_slogic(117),
    to_slogic(119),
    to_slogic(133),
    to_slogic(137),
    to_slogic(133),
    to_slogic(128),
    to_slogic(128),
    to_slogic(117),
    to_slogic(109),
    to_slogic(110),
    to_slogic(141),
    to_slogic(155),
    to_slogic(177),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(166),
    to_slogic(162),
    to_slogic(167),
    to_slogic(185),
    to_slogic(182),
    to_slogic(167),
    to_slogic(172),
    to_slogic(182),
    to_slogic(177),
    to_slogic(182),
    to_slogic(182),
    to_slogic(185),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(200),
    to_slogic(185),
    to_slogic(196),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(185),
    to_slogic(196),
    to_slogic(197),
    to_slogic(205),
    to_slogic(211),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(196),
    to_slogic(204),
    to_slogic(208),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(208),
    to_slogic(208),
    to_slogic(220),
    to_slogic(226),
    to_slogic(226),
    to_slogic(165),
    to_slogic(82),
    to_slogic(92),
    to_slogic(121),
    to_slogic(139),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(146),
    to_slogic(144),
    to_slogic(117),
    to_slogic(102),
    to_slogic(70),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(68),
    to_slogic(153),
    to_slogic(205),
    to_slogic(213),
    to_slogic(189),
    to_slogic(170),
    to_slogic(208),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(226),
    to_slogic(226),
    to_slogic(143),
    to_slogic(42),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(75),
    to_slogic(113),
    to_slogic(144),
    to_slogic(149),
    to_slogic(151),
    to_slogic(141),
    to_slogic(141),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(158),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(100),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(89),
    to_slogic(109),
    to_slogic(121),
    to_slogic(143),
    to_slogic(151),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(89),
    to_slogic(75),
    to_slogic(70),
    to_slogic(75),
    to_slogic(76),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(94),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(117),
    to_slogic(109),
    to_slogic(102),
    to_slogic(162),
    to_slogic(207),
    to_slogic(176),
    to_slogic(135),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(128),
    to_slogic(119),
    to_slogic(119),
    to_slogic(119),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(126),
    to_slogic(128),
    to_slogic(118),
    to_slogic(116),
    to_slogic(109),
    to_slogic(101),
    to_slogic(151),
    to_slogic(167),
    to_slogic(172),
    to_slogic(176),
    to_slogic(182),
    to_slogic(167),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(176),
    to_slogic(171),
    to_slogic(169),
    to_slogic(182),
    to_slogic(185),
    to_slogic(182),
    to_slogic(176),
    to_slogic(167),
    to_slogic(189),
    to_slogic(195),
    to_slogic(191),
    to_slogic(185),
    to_slogic(189),
    to_slogic(185),
    to_slogic(191),
    to_slogic(185),
    to_slogic(200),
    to_slogic(191),
    to_slogic(189),
    to_slogic(185),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(197),
    to_slogic(205),
    to_slogic(208),
    to_slogic(205),
    to_slogic(208),
    to_slogic(208),
    to_slogic(208),
    to_slogic(208),
    to_slogic(208),
    to_slogic(214),
    to_slogic(220),
    to_slogic(226),
    to_slogic(208),
    to_slogic(119),
    to_slogic(92),
    to_slogic(116),
    to_slogic(135),
    to_slogic(144),
    to_slogic(155),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(139),
    to_slogic(116),
    to_slogic(92),
    to_slogic(62),
    to_slogic(33),
    to_slogic(40),
    to_slogic(40),
    to_slogic(95),
    to_slogic(170),
    to_slogic(208),
    to_slogic(204),
    to_slogic(176),
    to_slogic(170),
    to_slogic(208),
    to_slogic(220),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(226),
    to_slogic(226),
    to_slogic(176),
    to_slogic(50),
    to_slogic(42),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(96),
    to_slogic(141),
    to_slogic(151),
    to_slogic(151),
    to_slogic(141),
    to_slogic(139),
    to_slogic(149),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(158),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(158),
    to_slogic(155),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(115),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(144),
    to_slogic(130),
    to_slogic(109),
    to_slogic(92),
    to_slogic(76),
    to_slogic(76),
    to_slogic(75),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(99),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(117),
    to_slogic(102),
    to_slogic(173),
    to_slogic(205),
    to_slogic(172),
    to_slogic(126),
    to_slogic(99),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(99),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(126),
    to_slogic(128),
    to_slogic(130),
    to_slogic(119),
    to_slogic(117),
    to_slogic(119),
    to_slogic(119),
    to_slogic(128),
    to_slogic(137),
    to_slogic(133),
    to_slogic(116),
    to_slogic(128),
    to_slogic(128),
    to_slogic(117),
    to_slogic(109),
    to_slogic(119),
    to_slogic(141),
    to_slogic(165),
    to_slogic(172),
    to_slogic(176),
    to_slogic(176),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(176),
    to_slogic(176),
    to_slogic(169),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(185),
    to_slogic(182),
    to_slogic(196),
    to_slogic(189),
    to_slogic(191),
    to_slogic(182),
    to_slogic(185),
    to_slogic(185),
    to_slogic(195),
    to_slogic(177),
    to_slogic(182),
    to_slogic(179),
    to_slogic(196),
    to_slogic(200),
    to_slogic(205),
    to_slogic(195),
    to_slogic(196),
    to_slogic(196),
    to_slogic(195),
    to_slogic(189),
    to_slogic(196),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(197),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(205),
    to_slogic(208),
    to_slogic(208),
    to_slogic(220),
    to_slogic(220),
    to_slogic(177),
    to_slogic(94),
    to_slogic(116),
    to_slogic(135),
    to_slogic(144),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(144),
    to_slogic(130),
    to_slogic(116),
    to_slogic(94),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(102),
    to_slogic(197),
    to_slogic(220),
    to_slogic(193),
    to_slogic(167),
    to_slogic(177),
    to_slogic(205),
    to_slogic(220),
    to_slogic(220),
    to_slogic(214),
    to_slogic(213),
    to_slogic(208),
    to_slogic(208),
    to_slogic(213),
    to_slogic(197),
    to_slogic(214),
    to_slogic(226),
    to_slogic(226),
    to_slogic(196),
    to_slogic(49),
    to_slogic(42),
    to_slogic(40),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(81),
    to_slogic(126),
    to_slogic(151),
    to_slogic(155),
    to_slogic(143),
    to_slogic(144),
    to_slogic(151),
    to_slogic(155),
    to_slogic(162),
    to_slogic(157),
    to_slogic(156),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(162),
    to_slogic(92),
    to_slogic(92),
    to_slogic(94),
    to_slogic(99),
    to_slogic(96),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(121),
    to_slogic(135),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(157),
    to_slogic(143),
    to_slogic(135),
    to_slogic(109),
    to_slogic(92),
    to_slogic(76),
    to_slogic(81),
    to_slogic(76),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(115),
    to_slogic(102),
    to_slogic(102),
    to_slogic(197),
    to_slogic(197),
    to_slogic(165),
    to_slogic(143),
    to_slogic(99),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(92),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(126),
    to_slogic(119),
    to_slogic(119),
    to_slogic(119),
    to_slogic(117),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(127),
    to_slogic(133),
    to_slogic(130),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(149),
    to_slogic(165),
    to_slogic(162),
    to_slogic(177),
    to_slogic(172),
    to_slogic(165),
    to_slogic(162),
    to_slogic(158),
    to_slogic(172),
    to_slogic(167),
    to_slogic(162),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(177),
    to_slogic(176),
    to_slogic(191),
    to_slogic(185),
    to_slogic(185),
    to_slogic(182),
    to_slogic(185),
    to_slogic(185),
    to_slogic(191),
    to_slogic(185),
    to_slogic(182),
    to_slogic(176),
    to_slogic(176),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(195),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(195),
    to_slogic(196),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(208),
    to_slogic(220),
    to_slogic(220),
    to_slogic(162),
    to_slogic(118),
    to_slogic(130),
    to_slogic(144),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(156),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(143),
    to_slogic(126),
    to_slogic(100),
    to_slogic(75),
    to_slogic(49),
    to_slogic(81),
    to_slogic(153),
    to_slogic(205),
    to_slogic(213),
    to_slogic(193),
    to_slogic(165),
    to_slogic(192),
    to_slogic(208),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(213),
    to_slogic(205),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(193),
    to_slogic(49),
    to_slogic(42),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(64),
    to_slogic(110),
    to_slogic(151),
    to_slogic(149),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(149),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(157),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(150),
    to_slogic(162),
    to_slogic(157),
    to_slogic(155),
    to_slogic(162),
    to_slogic(158),
    to_slogic(92),
    to_slogic(99),
    to_slogic(94),
    to_slogic(94),
    to_slogic(99),
    to_slogic(96),
    to_slogic(97),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(89),
    to_slogic(109),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(144),
    to_slogic(130),
    to_slogic(115),
    to_slogic(92),
    to_slogic(82),
    to_slogic(75),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(102),
    to_slogic(117),
    to_slogic(207),
    to_slogic(197),
    to_slogic(156),
    to_slogic(121),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(99),
    to_slogic(96),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(117),
    to_slogic(128),
    to_slogic(126),
    to_slogic(117),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(117),
    to_slogic(102),
    to_slogic(119),
    to_slogic(151),
    to_slogic(151),
    to_slogic(173),
    to_slogic(165),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(172),
    to_slogic(172),
    to_slogic(149),
    to_slogic(165),
    to_slogic(177),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(177),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(185),
    to_slogic(182),
    to_slogic(185),
    to_slogic(176),
    to_slogic(185),
    to_slogic(182),
    to_slogic(182),
    to_slogic(165),
    to_slogic(176),
    to_slogic(185),
    to_slogic(191),
    to_slogic(182),
    to_slogic(189),
    to_slogic(195),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(191),
    to_slogic(195),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(196),
    to_slogic(189),
    to_slogic(182),
    to_slogic(177),
    to_slogic(197),
    to_slogic(204),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(197),
    to_slogic(205),
    to_slogic(205),
    to_slogic(208),
    to_slogic(208),
    to_slogic(208),
    to_slogic(214),
    to_slogic(214),
    to_slogic(181),
    to_slogic(144),
    to_slogic(143),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(156),
    to_slogic(151),
    to_slogic(151),
    to_slogic(144),
    to_slogic(143),
    to_slogic(126),
    to_slogic(89),
    to_slogic(82),
    to_slogic(119),
    to_slogic(181),
    to_slogic(214),
    to_slogic(196),
    to_slogic(176),
    to_slogic(177),
    to_slogic(205),
    to_slogic(214),
    to_slogic(220),
    to_slogic(213),
    to_slogic(208),
    to_slogic(205),
    to_slogic(205),
    to_slogic(196),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(214),
    to_slogic(214),
    to_slogic(226),
    to_slogic(226),
    to_slogic(177),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(36),
    to_slogic(46),
    to_slogic(87),
    to_slogic(133),
    to_slogic(151),
    to_slogic(151),
    to_slogic(141),
    to_slogic(144),
    to_slogic(151),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(156),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(97),
    to_slogic(100),
    to_slogic(109),
    to_slogic(121),
    to_slogic(143),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(130),
    to_slogic(116),
    to_slogic(89),
    to_slogic(81),
    to_slogic(76),
    to_slogic(81),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(115),
    to_slogic(102),
    to_slogic(128),
    to_slogic(213),
    to_slogic(197),
    to_slogic(143),
    to_slogic(121),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(115),
    to_slogic(118),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(117),
    to_slogic(116),
    to_slogic(109),
    to_slogic(126),
    to_slogic(117),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(119),
    to_slogic(128),
    to_slogic(117),
    to_slogic(102),
    to_slogic(119),
    to_slogic(151),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(151),
    to_slogic(151),
    to_slogic(172),
    to_slogic(165),
    to_slogic(155),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(189),
    to_slogic(185),
    to_slogic(172),
    to_slogic(176),
    to_slogic(182),
    to_slogic(185),
    to_slogic(176),
    to_slogic(177),
    to_slogic(182),
    to_slogic(176),
    to_slogic(158),
    to_slogic(176),
    to_slogic(182),
    to_slogic(185),
    to_slogic(191),
    to_slogic(185),
    to_slogic(182),
    to_slogic(189),
    to_slogic(191),
    to_slogic(200),
    to_slogic(196),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(162),
    to_slogic(170),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(197),
    to_slogic(205),
    to_slogic(204),
    to_slogic(197),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(196),
    to_slogic(205),
    to_slogic(208),
    to_slogic(208),
    to_slogic(214),
    to_slogic(220),
    to_slogic(177),
    to_slogic(144),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(143),
    to_slogic(135),
    to_slogic(117),
    to_slogic(110),
    to_slogic(166),
    to_slogic(208),
    to_slogic(213),
    to_slogic(189),
    to_slogic(189),
    to_slogic(191),
    to_slogic(205),
    to_slogic(214),
    to_slogic(208),
    to_slogic(208),
    to_slogic(204),
    to_slogic(213),
    to_slogic(205),
    to_slogic(204),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(208),
    to_slogic(214),
    to_slogic(220),
    to_slogic(226),
    to_slogic(220),
    to_slogic(170),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(33),
    to_slogic(36),
    to_slogic(63),
    to_slogic(121),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(150),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(100),
    to_slogic(96),
    to_slogic(94),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(96),
    to_slogic(100),
    to_slogic(92),
    to_slogic(99),
    to_slogic(97),
    to_slogic(109),
    to_slogic(130),
    to_slogic(135),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(144),
    to_slogic(135),
    to_slogic(116),
    to_slogic(89),
    to_slogic(81),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(97),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(102),
    to_slogic(102),
    to_slogic(152),
    to_slogic(213),
    to_slogic(184),
    to_slogic(135),
    to_slogic(116),
    to_slogic(109),
    to_slogic(92),
    to_slogic(99),
    to_slogic(102),
    to_slogic(115),
    to_slogic(115),
    to_slogic(102),
    to_slogic(109),
    to_slogic(115),
    to_slogic(99),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(124),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(119),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(101),
    to_slogic(120),
    to_slogic(151),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(146),
    to_slogic(139),
    to_slogic(149),
    to_slogic(162),
    to_slogic(141),
    to_slogic(149),
    to_slogic(167),
    to_slogic(176),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(176),
    to_slogic(182),
    to_slogic(172),
    to_slogic(182),
    to_slogic(176),
    to_slogic(172),
    to_slogic(182),
    to_slogic(176),
    to_slogic(185),
    to_slogic(182),
    to_slogic(165),
    to_slogic(158),
    to_slogic(185),
    to_slogic(185),
    to_slogic(182),
    to_slogic(176),
    to_slogic(189),
    to_slogic(189),
    to_slogic(185),
    to_slogic(185),
    to_slogic(191),
    to_slogic(191),
    to_slogic(193),
    to_slogic(191),
    to_slogic(191),
    to_slogic(205),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(191),
    to_slogic(158),
    to_slogic(170),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(197),
    to_slogic(204),
    to_slogic(197),
    to_slogic(204),
    to_slogic(197),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(208),
    to_slogic(208),
    to_slogic(213),
    to_slogic(172),
    to_slogic(143),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(165),
    to_slogic(197),
    to_slogic(213),
    to_slogic(196),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(208),
    to_slogic(214),
    to_slogic(205),
    to_slogic(213),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(197),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(143),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(33),
    to_slogic(46),
    to_slogic(101),
    to_slogic(141),
    to_slogic(155),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(150),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(157),
    to_slogic(149),
    to_slogic(155),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(130),
    to_slogic(121),
    to_slogic(89),
    to_slogic(81),
    to_slogic(81),
    to_slogic(81),
    to_slogic(89),
    to_slogic(82),
    to_slogic(100),
    to_slogic(99),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(100),
    to_slogic(99),
    to_slogic(173),
    to_slogic(207),
    to_slogic(165),
    to_slogic(135),
    to_slogic(126),
    to_slogic(116),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(99),
    to_slogic(102),
    to_slogic(99),
    to_slogic(102),
    to_slogic(121),
    to_slogic(117),
    to_slogic(118),
    to_slogic(109),
    to_slogic(124),
    to_slogic(128),
    to_slogic(128),
    to_slogic(124),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(109),
    to_slogic(127),
    to_slogic(144),
    to_slogic(155),
    to_slogic(162),
    to_slogic(151),
    to_slogic(152),
    to_slogic(149),
    to_slogic(151),
    to_slogic(151),
    to_slogic(139),
    to_slogic(151),
    to_slogic(162),
    to_slogic(165),
    to_slogic(172),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(167),
    to_slogic(172),
    to_slogic(172),
    to_slogic(182),
    to_slogic(185),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(165),
    to_slogic(172),
    to_slogic(176),
    to_slogic(176),
    to_slogic(185),
    to_slogic(185),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(189),
    to_slogic(185),
    to_slogic(182),
    to_slogic(185),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(182),
    to_slogic(170),
    to_slogic(176),
    to_slogic(189),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(197),
    to_slogic(204),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(197),
    to_slogic(208),
    to_slogic(205),
    to_slogic(191),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(162),
    to_slogic(200),
    to_slogic(214),
    to_slogic(207),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(197),
    to_slogic(208),
    to_slogic(208),
    to_slogic(213),
    to_slogic(205),
    to_slogic(204),
    to_slogic(197),
    to_slogic(196),
    to_slogic(197),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(114),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(46),
    to_slogic(81),
    to_slogic(127),
    to_slogic(151),
    to_slogic(149),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(157),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(155),
    to_slogic(150),
    to_slogic(157),
    to_slogic(155),
    to_slogic(96),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(94),
    to_slogic(97),
    to_slogic(109),
    to_slogic(115),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(152),
    to_slogic(161),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(156),
    to_slogic(151),
    to_slogic(135),
    to_slogic(116),
    to_slogic(97),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(99),
    to_slogic(102),
    to_slogic(183),
    to_slogic(205),
    to_slogic(165),
    to_slogic(143),
    to_slogic(121),
    to_slogic(116),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(117),
    to_slogic(117),
    to_slogic(119),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(126),
    to_slogic(109),
    to_slogic(117),
    to_slogic(134),
    to_slogic(143),
    to_slogic(149),
    to_slogic(152),
    to_slogic(150),
    to_slogic(146),
    to_slogic(146),
    to_slogic(155),
    to_slogic(155),
    to_slogic(125),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(155),
    to_slogic(172),
    to_slogic(182),
    to_slogic(176),
    to_slogic(162),
    to_slogic(165),
    to_slogic(167),
    to_slogic(162),
    to_slogic(167),
    to_slogic(185),
    to_slogic(182),
    to_slogic(185),
    to_slogic(165),
    to_slogic(155),
    to_slogic(172),
    to_slogic(182),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(185),
    to_slogic(176),
    to_slogic(182),
    to_slogic(196),
    to_slogic(200),
    to_slogic(182),
    to_slogic(189),
    to_slogic(179),
    to_slogic(165),
    to_slogic(191),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(185),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(196),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(181),
    to_slogic(196),
    to_slogic(191),
    to_slogic(196),
    to_slogic(197),
    to_slogic(205),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(144),
    to_slogic(155),
    to_slogic(182),
    to_slogic(205),
    to_slogic(204),
    to_slogic(189),
    to_slogic(193),
    to_slogic(176),
    to_slogic(191),
    to_slogic(205),
    to_slogic(213),
    to_slogic(208),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(81),
    to_slogic(49),
    to_slogic(50),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(69),
    to_slogic(109),
    to_slogic(141),
    to_slogic(155),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(100),
    to_slogic(102),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(97),
    to_slogic(97),
    to_slogic(100),
    to_slogic(109),
    to_slogic(130),
    to_slogic(143),
    to_slogic(152),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(109),
    to_slogic(97),
    to_slogic(75),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(99),
    to_slogic(102),
    to_slogic(207),
    to_slogic(197),
    to_slogic(172),
    to_slogic(143),
    to_slogic(130),
    to_slogic(116),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(126),
    to_slogic(117),
    to_slogic(109),
    to_slogic(128),
    to_slogic(119),
    to_slogic(117),
    to_slogic(119),
    to_slogic(134),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(144),
    to_slogic(146),
    to_slogic(139),
    to_slogic(155),
    to_slogic(137),
    to_slogic(127),
    to_slogic(151),
    to_slogic(155),
    to_slogic(155),
    to_slogic(165),
    to_slogic(172),
    to_slogic(158),
    to_slogic(172),
    to_slogic(172),
    to_slogic(167),
    to_slogic(172),
    to_slogic(165),
    to_slogic(176),
    to_slogic(172),
    to_slogic(167),
    to_slogic(176),
    to_slogic(166),
    to_slogic(157),
    to_slogic(167),
    to_slogic(182),
    to_slogic(176),
    to_slogic(176),
    to_slogic(172),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(185),
    to_slogic(172),
    to_slogic(182),
    to_slogic(185),
    to_slogic(185),
    to_slogic(185),
    to_slogic(167),
    to_slogic(162),
    to_slogic(176),
    to_slogic(182),
    to_slogic(185),
    to_slogic(189),
    to_slogic(176),
    to_slogic(176),
    to_slogic(185),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(196),
    to_slogic(185),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(177),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(204),
    to_slogic(170),
    to_slogic(144),
    to_slogic(155),
    to_slogic(179),
    to_slogic(204),
    to_slogic(204),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(189),
    to_slogic(196),
    to_slogic(214),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(196),
    to_slogic(205),
    to_slogic(197),
    to_slogic(205),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(226),
    to_slogic(204),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(69),
    to_slogic(96),
    to_slogic(133),
    to_slogic(151),
    to_slogic(144),
    to_slogic(141),
    to_slogic(151),
    to_slogic(149),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(100),
    to_slogic(96),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(97),
    to_slogic(109),
    to_slogic(115),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(161),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(116),
    to_slogic(99),
    to_slogic(81),
    to_slogic(76),
    to_slogic(81),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(96),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(99),
    to_slogic(92),
    to_slogic(117),
    to_slogic(213),
    to_slogic(196),
    to_slogic(165),
    to_slogic(151),
    to_slogic(130),
    to_slogic(116),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(118),
    to_slogic(109),
    to_slogic(124),
    to_slogic(109),
    to_slogic(117),
    to_slogic(126),
    to_slogic(128),
    to_slogic(124),
    to_slogic(110),
    to_slogic(133),
    to_slogic(139),
    to_slogic(146),
    to_slogic(155),
    to_slogic(151),
    to_slogic(137),
    to_slogic(139),
    to_slogic(155),
    to_slogic(137),
    to_slogic(125),
    to_slogic(151),
    to_slogic(151),
    to_slogic(165),
    to_slogic(155),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(157),
    to_slogic(162),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(167),
    to_slogic(176),
    to_slogic(165),
    to_slogic(156),
    to_slogic(157),
    to_slogic(171),
    to_slogic(176),
    to_slogic(167),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(172),
    to_slogic(176),
    to_slogic(176),
    to_slogic(172),
    to_slogic(182),
    to_slogic(176),
    to_slogic(185),
    to_slogic(185),
    to_slogic(191),
    to_slogic(189),
    to_slogic(176),
    to_slogic(172),
    to_slogic(182),
    to_slogic(185),
    to_slogic(185),
    to_slogic(189),
    to_slogic(177),
    to_slogic(176),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(189),
    to_slogic(191),
    to_slogic(185),
    to_slogic(177),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(185),
    to_slogic(177),
    to_slogic(191),
    to_slogic(191),
    to_slogic(181),
    to_slogic(191),
    to_slogic(196),
    to_slogic(172),
    to_slogic(189),
    to_slogic(204),
    to_slogic(207),
    to_slogic(176),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(197),
    to_slogic(204),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(214),
    to_slogic(205),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(189),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(69),
    to_slogic(81),
    to_slogic(117),
    to_slogic(141),
    to_slogic(151),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(157),
    to_slogic(162),
    to_slogic(155),
    to_slogic(157),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(102),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(157),
    to_slogic(151),
    to_slogic(130),
    to_slogic(121),
    to_slogic(89),
    to_slogic(81),
    to_slogic(81),
    to_slogic(76),
    to_slogic(89),
    to_slogic(89),
    to_slogic(92),
    to_slogic(89),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(137),
    to_slogic(213),
    to_slogic(191),
    to_slogic(172),
    to_slogic(151),
    to_slogic(144),
    to_slogic(121),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(115),
    to_slogic(109),
    to_slogic(115),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(119),
    to_slogic(124),
    to_slogic(128),
    to_slogic(117),
    to_slogic(109),
    to_slogic(128),
    to_slogic(151),
    to_slogic(149),
    to_slogic(151),
    to_slogic(146),
    to_slogic(137),
    to_slogic(146),
    to_slogic(143),
    to_slogic(128),
    to_slogic(133),
    to_slogic(141),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(172),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(172),
    to_slogic(182),
    to_slogic(182),
    to_slogic(171),
    to_slogic(162),
    to_slogic(155),
    to_slogic(165),
    to_slogic(182),
    to_slogic(176),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(167),
    to_slogic(182),
    to_slogic(167),
    to_slogic(176),
    to_slogic(167),
    to_slogic(167),
    to_slogic(176),
    to_slogic(176),
    to_slogic(185),
    to_slogic(191),
    to_slogic(182),
    to_slogic(176),
    to_slogic(177),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(177),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(179),
    to_slogic(176),
    to_slogic(185),
    to_slogic(185),
    to_slogic(185),
    to_slogic(185),
    to_slogic(177),
    to_slogic(185),
    to_slogic(185),
    to_slogic(177),
    to_slogic(176),
    to_slogic(181),
    to_slogic(185),
    to_slogic(189),
    to_slogic(196),
    to_slogic(193),
    to_slogic(207),
    to_slogic(189),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(197),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(220),
    to_slogic(153),
    to_slogic(40),
    to_slogic(40),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(75),
    to_slogic(101),
    to_slogic(141),
    to_slogic(151),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(155),
    to_slogic(157),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(102),
    to_slogic(96),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(97),
    to_slogic(100),
    to_slogic(116),
    to_slogic(121),
    to_slogic(143),
    to_slogic(151),
    to_slogic(161),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(89),
    to_slogic(76),
    to_slogic(70),
    to_slogic(81),
    to_slogic(92),
    to_slogic(89),
    to_slogic(99),
    to_slogic(94),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(115),
    to_slogic(100),
    to_slogic(99),
    to_slogic(102),
    to_slogic(92),
    to_slogic(157),
    to_slogic(213),
    to_slogic(191),
    to_slogic(184),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(121),
    to_slogic(126),
    to_slogic(109),
    to_slogic(109),
    to_slogic(118),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(117),
    to_slogic(100),
    to_slogic(109),
    to_slogic(124),
    to_slogic(117),
    to_slogic(126),
    to_slogic(124),
    to_slogic(110),
    to_slogic(119),
    to_slogic(146),
    to_slogic(141),
    to_slogic(152),
    to_slogic(137),
    to_slogic(133),
    to_slogic(146),
    to_slogic(149),
    to_slogic(133),
    to_slogic(133),
    to_slogic(141),
    to_slogic(146),
    to_slogic(151),
    to_slogic(151),
    to_slogic(155),
    to_slogic(139),
    to_slogic(155),
    to_slogic(149),
    to_slogic(162),
    to_slogic(172),
    to_slogic(176),
    to_slogic(165),
    to_slogic(165),
    to_slogic(167),
    to_slogic(165),
    to_slogic(149),
    to_slogic(172),
    to_slogic(167),
    to_slogic(177),
    to_slogic(176),
    to_slogic(167),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(172),
    to_slogic(167),
    to_slogic(172),
    to_slogic(182),
    to_slogic(172),
    to_slogic(176),
    to_slogic(185),
    to_slogic(185),
    to_slogic(182),
    to_slogic(182),
    to_slogic(179),
    to_slogic(176),
    to_slogic(185),
    to_slogic(185),
    to_slogic(191),
    to_slogic(191),
    to_slogic(185),
    to_slogic(189),
    to_slogic(191),
    to_slogic(185),
    to_slogic(176),
    to_slogic(182),
    to_slogic(172),
    to_slogic(176),
    to_slogic(185),
    to_slogic(181),
    to_slogic(185),
    to_slogic(182),
    to_slogic(179),
    to_slogic(177),
    to_slogic(165),
    to_slogic(165),
    to_slogic(170),
    to_slogic(189),
    to_slogic(196),
    to_slogic(193),
    to_slogic(182),
    to_slogic(170),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(214),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(205),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(189),
    to_slogic(182),
    to_slogic(191),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(220),
    to_slogic(213),
    to_slogic(102),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(46),
    to_slogic(64),
    to_slogic(96),
    to_slogic(126),
    to_slogic(151),
    to_slogic(151),
    to_slogic(143),
    to_slogic(141),
    to_slogic(151),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(150),
    to_slogic(162),
    to_slogic(150),
    to_slogic(94),
    to_slogic(99),
    to_slogic(99),
    to_slogic(96),
    to_slogic(102),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(165),
    to_slogic(165),
    to_slogic(151),
    to_slogic(130),
    to_slogic(121),
    to_slogic(99),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(81),
    to_slogic(92),
    to_slogic(97),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(97),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(82),
    to_slogic(165),
    to_slogic(213),
    to_slogic(183),
    to_slogic(176),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(116),
    to_slogic(100),
    to_slogic(102),
    to_slogic(118),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(126),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(110),
    to_slogic(128),
    to_slogic(134),
    to_slogic(137),
    to_slogic(149),
    to_slogic(146),
    to_slogic(139),
    to_slogic(146),
    to_slogic(143),
    to_slogic(128),
    to_slogic(120),
    to_slogic(146),
    to_slogic(155),
    to_slogic(152),
    to_slogic(151),
    to_slogic(155),
    to_slogic(139),
    to_slogic(146),
    to_slogic(139),
    to_slogic(155),
    to_slogic(165),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(165),
    to_slogic(139),
    to_slogic(162),
    to_slogic(176),
    to_slogic(176),
    to_slogic(172),
    to_slogic(162),
    to_slogic(162),
    to_slogic(176),
    to_slogic(172),
    to_slogic(177),
    to_slogic(182),
    to_slogic(176),
    to_slogic(167),
    to_slogic(176),
    to_slogic(176),
    to_slogic(172),
    to_slogic(172),
    to_slogic(167),
    to_slogic(172),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(177),
    to_slogic(182),
    to_slogic(177),
    to_slogic(176),
    to_slogic(185),
    to_slogic(191),
    to_slogic(191),
    to_slogic(185),
    to_slogic(185),
    to_slogic(179),
    to_slogic(185),
    to_slogic(185),
    to_slogic(170),
    to_slogic(176),
    to_slogic(170),
    to_slogic(176),
    to_slogic(177),
    to_slogic(185),
    to_slogic(165),
    to_slogic(170),
    to_slogic(167),
    to_slogic(162),
    to_slogic(176),
    to_slogic(196),
    to_slogic(193),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(196),
    to_slogic(197),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(205),
    to_slogic(205),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(196),
    to_slogic(176),
    to_slogic(165),
    to_slogic(182),
    to_slogic(196),
    to_slogic(205),
    to_slogic(204),
    to_slogic(214),
    to_slogic(214),
    to_slogic(207),
    to_slogic(68),
    to_slogic(36),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(44),
    to_slogic(63),
    to_slogic(110),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(150),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(99),
    to_slogic(100),
    to_slogic(96),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(94),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(161),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(92),
    to_slogic(82),
    to_slogic(81),
    to_slogic(81),
    to_slogic(92),
    to_slogic(99),
    to_slogic(89),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(173),
    to_slogic(213),
    to_slogic(184),
    to_slogic(172),
    to_slogic(165),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(130),
    to_slogic(121),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(118),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(102),
    to_slogic(102),
    to_slogic(128),
    to_slogic(146),
    to_slogic(137),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(144),
    to_slogic(143),
    to_slogic(119),
    to_slogic(128),
    to_slogic(146),
    to_slogic(152),
    to_slogic(139),
    to_slogic(155),
    to_slogic(155),
    to_slogic(151),
    to_slogic(133),
    to_slogic(141),
    to_slogic(151),
    to_slogic(151),
    to_slogic(162),
    to_slogic(155),
    to_slogic(167),
    to_slogic(165),
    to_slogic(151),
    to_slogic(157),
    to_slogic(172),
    to_slogic(176),
    to_slogic(176),
    to_slogic(172),
    to_slogic(167),
    to_slogic(165),
    to_slogic(166),
    to_slogic(176),
    to_slogic(172),
    to_slogic(177),
    to_slogic(176),
    to_slogic(172),
    to_slogic(157),
    to_slogic(162),
    to_slogic(167),
    to_slogic(172),
    to_slogic(156),
    to_slogic(172),
    to_slogic(176),
    to_slogic(167),
    to_slogic(176),
    to_slogic(167),
    to_slogic(176),
    to_slogic(182),
    to_slogic(185),
    to_slogic(185),
    to_slogic(177),
    to_slogic(182),
    to_slogic(185),
    to_slogic(189),
    to_slogic(185),
    to_slogic(177),
    to_slogic(176),
    to_slogic(179),
    to_slogic(177),
    to_slogic(185),
    to_slogic(179),
    to_slogic(172),
    to_slogic(172),
    to_slogic(182),
    to_slogic(170),
    to_slogic(167),
    to_slogic(162),
    to_slogic(165),
    to_slogic(191),
    to_slogic(207),
    to_slogic(189),
    to_slogic(176),
    to_slogic(185),
    to_slogic(191),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(196),
    to_slogic(204),
    to_slogic(197),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(176),
    to_slogic(162),
    to_slogic(156),
    to_slogic(176),
    to_slogic(191),
    to_slogic(193),
    to_slogic(189),
    to_slogic(205),
    to_slogic(213),
    to_slogic(153),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(81),
    to_slogic(125),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(144),
    to_slogic(157),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(150),
    to_slogic(162),
    to_slogic(150),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(162),
    to_slogic(157),
    to_slogic(155),
    to_slogic(99),
    to_slogic(94),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(130),
    to_slogic(144),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(165),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(92),
    to_slogic(81),
    to_slogic(76),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(94),
    to_slogic(99),
    to_slogic(99),
    to_slogic(96),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(97),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(173),
    to_slogic(207),
    to_slogic(184),
    to_slogic(172),
    to_slogic(156),
    to_slogic(161),
    to_slogic(135),
    to_slogic(143),
    to_slogic(135),
    to_slogic(130),
    to_slogic(116),
    to_slogic(109),
    to_slogic(99),
    to_slogic(89),
    to_slogic(109),
    to_slogic(102),
    to_slogic(117),
    to_slogic(124),
    to_slogic(109),
    to_slogic(102),
    to_slogic(119),
    to_slogic(139),
    to_slogic(146),
    to_slogic(133),
    to_slogic(134),
    to_slogic(144),
    to_slogic(146),
    to_slogic(139),
    to_slogic(119),
    to_slogic(119),
    to_slogic(146),
    to_slogic(141),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(141),
    to_slogic(141),
    to_slogic(165),
    to_slogic(151),
    to_slogic(141),
    to_slogic(165),
    to_slogic(176),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(167),
    to_slogic(167),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(172),
    to_slogic(172),
    to_slogic(162),
    to_slogic(165),
    to_slogic(167),
    to_slogic(165),
    to_slogic(162),
    to_slogic(167),
    to_slogic(172),
    to_slogic(167),
    to_slogic(162),
    to_slogic(162),
    to_slogic(172),
    to_slogic(172),
    to_slogic(167),
    to_slogic(176),
    to_slogic(176),
    to_slogic(185),
    to_slogic(185),
    to_slogic(179),
    to_slogic(182),
    to_slogic(179),
    to_slogic(176),
    to_slogic(176),
    to_slogic(165),
    to_slogic(176),
    to_slogic(179),
    to_slogic(185),
    to_slogic(177),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(167),
    to_slogic(176),
    to_slogic(193),
    to_slogic(193),
    to_slogic(182),
    to_slogic(189),
    to_slogic(191),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(193),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(205),
    to_slogic(204),
    to_slogic(197),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(189),
    to_slogic(156),
    to_slogic(158),
    to_slogic(157),
    to_slogic(182),
    to_slogic(166),
    to_slogic(158),
    to_slogic(185),
    to_slogic(204),
    to_slogic(213),
    to_slogic(91),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(50),
    to_slogic(75),
    to_slogic(75),
    to_slogic(117),
    to_slogic(141),
    to_slogic(155),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(157),
    to_slogic(162),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(155),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(92),
    to_slogic(94),
    to_slogic(92),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(135),
    to_slogic(143),
    to_slogic(157),
    to_slogic(161),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(151),
    to_slogic(135),
    to_slogic(116),
    to_slogic(92),
    to_slogic(81),
    to_slogic(75),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(96),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(87),
    to_slogic(178),
    to_slogic(197),
    to_slogic(183),
    to_slogic(169),
    to_slogic(165),
    to_slogic(157),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(135),
    to_slogic(121),
    to_slogic(115),
    to_slogic(102),
    to_slogic(99),
    to_slogic(89),
    to_slogic(115),
    to_slogic(116),
    to_slogic(109),
    to_slogic(102),
    to_slogic(128),
    to_slogic(146),
    to_slogic(133),
    to_slogic(146),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(139),
    to_slogic(119),
    to_slogic(119),
    to_slogic(133),
    to_slogic(146),
    to_slogic(152),
    to_slogic(151),
    to_slogic(146),
    to_slogic(137),
    to_slogic(141),
    to_slogic(151),
    to_slogic(155),
    to_slogic(141),
    to_slogic(144),
    to_slogic(151),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(155),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(167),
    to_slogic(169),
    to_slogic(155),
    to_slogic(166),
    to_slogic(172),
    to_slogic(157),
    to_slogic(165),
    to_slogic(166),
    to_slogic(172),
    to_slogic(157),
    to_slogic(165),
    to_slogic(155),
    to_slogic(158),
    to_slogic(165),
    to_slogic(165),
    to_slogic(176),
    to_slogic(176),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(185),
    to_slogic(177),
    to_slogic(170),
    to_slogic(172),
    to_slogic(170),
    to_slogic(176),
    to_slogic(172),
    to_slogic(162),
    to_slogic(165),
    to_slogic(185),
    to_slogic(176),
    to_slogic(162),
    to_slogic(156),
    to_slogic(149),
    to_slogic(182),
    to_slogic(193),
    to_slogic(198),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(196),
    to_slogic(167),
    to_slogic(155),
    to_slogic(158),
    to_slogic(176),
    to_slogic(166),
    to_slogic(134),
    to_slogic(156),
    to_slogic(185),
    to_slogic(207),
    to_slogic(177),
    to_slogic(49),
    to_slogic(42),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(50),
    to_slogic(64),
    to_slogic(81),
    to_slogic(101),
    to_slogic(133),
    to_slogic(151),
    to_slogic(151),
    to_slogic(139),
    to_slogic(141),
    to_slogic(157),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(150),
    to_slogic(156),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(92),
    to_slogic(94),
    to_slogic(92),
    to_slogic(89),
    to_slogic(100),
    to_slogic(99),
    to_slogic(115),
    to_slogic(130),
    to_slogic(144),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(99),
    to_slogic(81),
    to_slogic(77),
    to_slogic(82),
    to_slogic(82),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(96),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(97),
    to_slogic(92),
    to_slogic(89),
    to_slogic(183),
    to_slogic(196),
    to_slogic(175),
    to_slogic(172),
    to_slogic(161),
    to_slogic(161),
    to_slogic(151),
    to_slogic(143),
    to_slogic(135),
    to_slogic(144),
    to_slogic(121),
    to_slogic(100),
    to_slogic(102),
    to_slogic(99),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(99),
    to_slogic(127),
    to_slogic(146),
    to_slogic(139),
    to_slogic(139),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(119),
    to_slogic(119),
    to_slogic(139),
    to_slogic(137),
    to_slogic(146),
    to_slogic(152),
    to_slogic(141),
    to_slogic(137),
    to_slogic(146),
    to_slogic(137),
    to_slogic(151),
    to_slogic(137),
    to_slogic(151),
    to_slogic(155),
    to_slogic(155),
    to_slogic(146),
    to_slogic(146),
    to_slogic(162),
    to_slogic(165),
    to_slogic(155),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(172),
    to_slogic(169),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(162),
    to_slogic(157),
    to_slogic(162),
    to_slogic(172),
    to_slogic(165),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(167),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(167),
    to_slogic(165),
    to_slogic(172),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(162),
    to_slogic(158),
    to_slogic(189),
    to_slogic(193),
    to_slogic(171),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(196),
    to_slogic(193),
    to_slogic(191),
    to_slogic(189),
    to_slogic(196),
    to_slogic(189),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(197),
    to_slogic(205),
    to_slogic(214),
    to_slogic(205),
    to_slogic(204),
    to_slogic(182),
    to_slogic(149),
    to_slogic(165),
    to_slogic(176),
    to_slogic(166),
    to_slogic(132),
    to_slogic(151),
    to_slogic(165),
    to_slogic(182),
    to_slogic(205),
    to_slogic(144),
    to_slogic(36),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(50),
    to_slogic(69),
    to_slogic(82),
    to_slogic(127),
    to_slogic(151),
    to_slogic(151),
    to_slogic(144),
    to_slogic(151),
    to_slogic(151),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(162),
    to_slogic(158),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(89),
    to_slogic(92),
    to_slogic(100),
    to_slogic(89),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(121),
    to_slogic(135),
    to_slogic(143),
    to_slogic(152),
    to_slogic(161),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(92),
    to_slogic(82),
    to_slogic(76),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(96),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(94),
    to_slogic(100),
    to_slogic(89),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(99),
    to_slogic(198),
    to_slogic(191),
    to_slogic(184),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(144),
    to_slogic(121),
    to_slogic(121),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(115),
    to_slogic(102),
    to_slogic(128),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(133),
    to_slogic(128),
    to_slogic(137),
    to_slogic(128),
    to_slogic(118),
    to_slogic(127),
    to_slogic(133),
    to_slogic(146),
    to_slogic(146),
    to_slogic(143),
    to_slogic(133),
    to_slogic(146),
    to_slogic(139),
    to_slogic(144),
    to_slogic(132),
    to_slogic(139),
    to_slogic(141),
    to_slogic(155),
    to_slogic(149),
    to_slogic(149),
    to_slogic(151),
    to_slogic(157),
    to_slogic(155),
    to_slogic(162),
    to_slogic(157),
    to_slogic(152),
    to_slogic(151),
    to_slogic(165),
    to_slogic(162),
    to_slogic(172),
    to_slogic(155),
    to_slogic(157),
    to_slogic(155),
    to_slogic(162),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(162),
    to_slogic(155),
    to_slogic(141),
    to_slogic(162),
    to_slogic(162),
    to_slogic(167),
    to_slogic(165),
    to_slogic(172),
    to_slogic(158),
    to_slogic(165),
    to_slogic(162),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(167),
    to_slogic(169),
    to_slogic(158),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(162),
    to_slogic(149),
    to_slogic(156),
    to_slogic(182),
    to_slogic(189),
    to_slogic(182),
    to_slogic(171),
    to_slogic(182),
    to_slogic(193),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(189),
    to_slogic(196),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(196),
    to_slogic(205),
    to_slogic(204),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(196),
    to_slogic(155),
    to_slogic(158),
    to_slogic(176),
    to_slogic(166),
    to_slogic(141),
    to_slogic(149),
    to_slogic(162),
    to_slogic(172),
    to_slogic(189),
    to_slogic(213),
    to_slogic(91),
    to_slogic(42),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(109),
    to_slogic(141),
    to_slogic(155),
    to_slogic(151),
    to_slogic(149),
    to_slogic(141),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(102),
    to_slogic(115),
    to_slogic(130),
    to_slogic(143),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(94),
    to_slogic(81),
    to_slogic(81),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(97),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(89),
    to_slogic(82),
    to_slogic(99),
    to_slogic(197),
    to_slogic(191),
    to_slogic(184),
    to_slogic(184),
    to_slogic(172),
    to_slogic(156),
    to_slogic(151),
    to_slogic(151),
    to_slogic(143),
    to_slogic(143),
    to_slogic(135),
    to_slogic(121),
    to_slogic(116),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(119),
    to_slogic(133),
    to_slogic(146),
    to_slogic(139),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(128),
    to_slogic(110),
    to_slogic(119),
    to_slogic(133),
    to_slogic(146),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(133),
    to_slogic(146),
    to_slogic(137),
    to_slogic(127),
    to_slogic(133),
    to_slogic(151),
    to_slogic(151),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(151),
    to_slogic(155),
    to_slogic(157),
    to_slogic(151),
    to_slogic(151),
    to_slogic(162),
    to_slogic(162),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(143),
    to_slogic(161),
    to_slogic(162),
    to_slogic(169),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(144),
    to_slogic(157),
    to_slogic(155),
    to_slogic(165),
    to_slogic(167),
    to_slogic(157),
    to_slogic(165),
    to_slogic(167),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(162),
    to_slogic(162),
    to_slogic(165),
    to_slogic(157),
    to_slogic(162),
    to_slogic(172),
    to_slogic(157),
    to_slogic(165),
    to_slogic(149),
    to_slogic(149),
    to_slogic(176),
    to_slogic(182),
    to_slogic(189),
    to_slogic(177),
    to_slogic(183),
    to_slogic(182),
    to_slogic(193),
    to_slogic(200),
    to_slogic(193),
    to_slogic(198),
    to_slogic(193),
    to_slogic(189),
    to_slogic(182),
    to_slogic(193),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(204),
    to_slogic(197),
    to_slogic(204),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(204),
    to_slogic(167),
    to_slogic(155),
    to_slogic(172),
    to_slogic(156),
    to_slogic(144),
    to_slogic(165),
    to_slogic(166),
    to_slogic(151),
    to_slogic(158),
    to_slogic(204),
    to_slogic(177),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(87),
    to_slogic(133),
    to_slogic(149),
    to_slogic(151),
    to_slogic(143),
    to_slogic(141),
    to_slogic(155),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(150),
    to_slogic(162),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(158),
    to_slogic(92),
    to_slogic(94),
    to_slogic(102),
    to_slogic(92),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(121),
    to_slogic(135),
    to_slogic(143),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(144),
    to_slogic(124),
    to_slogic(102),
    to_slogic(76),
    to_slogic(76),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(97),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(89),
    to_slogic(109),
    to_slogic(207),
    to_slogic(191),
    to_slogic(197),
    to_slogic(176),
    to_slogic(176),
    to_slogic(165),
    to_slogic(161),
    to_slogic(151),
    to_slogic(143),
    to_slogic(143),
    to_slogic(135),
    to_slogic(130),
    to_slogic(115),
    to_slogic(99),
    to_slogic(92),
    to_slogic(119),
    to_slogic(144),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(128),
    to_slogic(137),
    to_slogic(128),
    to_slogic(119),
    to_slogic(119),
    to_slogic(133),
    to_slogic(146),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(146),
    to_slogic(125),
    to_slogic(119),
    to_slogic(134),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(134),
    to_slogic(146),
    to_slogic(155),
    to_slogic(157),
    to_slogic(155),
    to_slogic(155),
    to_slogic(157),
    to_slogic(151),
    to_slogic(154),
    to_slogic(162),
    to_slogic(155),
    to_slogic(160),
    to_slogic(148),
    to_slogic(143),
    to_slogic(134),
    to_slogic(126),
    to_slogic(125),
    to_slogic(127),
    to_slogic(143),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(162),
    to_slogic(162),
    to_slogic(157),
    to_slogic(162),
    to_slogic(172),
    to_slogic(155),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(167),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(151),
    to_slogic(158),
    to_slogic(149),
    to_slogic(149),
    to_slogic(167),
    to_slogic(182),
    to_slogic(189),
    to_slogic(177),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(204),
    to_slogic(204),
    to_slogic(193),
    to_slogic(189),
    to_slogic(176),
    to_slogic(189),
    to_slogic(176),
    to_slogic(191),
    to_slogic(189),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(214),
    to_slogic(205),
    to_slogic(214),
    to_slogic(191),
    to_slogic(149),
    to_slogic(167),
    to_slogic(156),
    to_slogic(149),
    to_slogic(162),
    to_slogic(137),
    to_slogic(119),
    to_slogic(141),
    to_slogic(177),
    to_slogic(220),
    to_slogic(132),
    to_slogic(40),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(69),
    to_slogic(101),
    to_slogic(141),
    to_slogic(151),
    to_slogic(151),
    to_slogic(149),
    to_slogic(151),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(158),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(162),
    to_slogic(150),
    to_slogic(99),
    to_slogic(100),
    to_slogic(92),
    to_slogic(102),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(115),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(161),
    to_slogic(152),
    to_slogic(143),
    to_slogic(121),
    to_slogic(92),
    to_slogic(81),
    to_slogic(70),
    to_slogic(76),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(100),
    to_slogic(97),
    to_slogic(100),
    to_slogic(97),
    to_slogic(99),
    to_slogic(89),
    to_slogic(82),
    to_slogic(100),
    to_slogic(207),
    to_slogic(205),
    to_slogic(191),
    to_slogic(191),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(143),
    to_slogic(143),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(92),
    to_slogic(102),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(127),
    to_slogic(139),
    to_slogic(128),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(146),
    to_slogic(139),
    to_slogic(133),
    to_slogic(146),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(127),
    to_slogic(134),
    to_slogic(133),
    to_slogic(151),
    to_slogic(151),
    to_slogic(133),
    to_slogic(134),
    to_slogic(149),
    to_slogic(155),
    to_slogic(162),
    to_slogic(151),
    to_slogic(141),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(155),
    to_slogic(144),
    to_slogic(126),
    to_slogic(142),
    to_slogic(144),
    to_slogic(133),
    to_slogic(96),
    to_slogic(101),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(165),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(149),
    to_slogic(157),
    to_slogic(157),
    to_slogic(155),
    to_slogic(165),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(155),
    to_slogic(167),
    to_slogic(193),
    to_slogic(182),
    to_slogic(177),
    to_slogic(171),
    to_slogic(185),
    to_slogic(200),
    to_slogic(193),
    to_slogic(204),
    to_slogic(193),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(197),
    to_slogic(204),
    to_slogic(205),
    to_slogic(197),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(208),
    to_slogic(205),
    to_slogic(158),
    to_slogic(165),
    to_slogic(155),
    to_slogic(149),
    to_slogic(118),
    to_slogic(107),
    to_slogic(96),
    to_slogic(127),
    to_slogic(158),
    to_slogic(204),
    to_slogic(213),
    to_slogic(68),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(81),
    to_slogic(134),
    to_slogic(149),
    to_slogic(151),
    to_slogic(151),
    to_slogic(141),
    to_slogic(149),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(150),
    to_slogic(162),
    to_slogic(150),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(102),
    to_slogic(92),
    to_slogic(100),
    to_slogic(94),
    to_slogic(92),
    to_slogic(102),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(121),
    to_slogic(130),
    to_slogic(143),
    to_slogic(157),
    to_slogic(156),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(135),
    to_slogic(116),
    to_slogic(97),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(99),
    to_slogic(96),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(89),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(89),
    to_slogic(97),
    to_slogic(81),
    to_slogic(100),
    to_slogic(207),
    to_slogic(197),
    to_slogic(197),
    to_slogic(183),
    to_slogic(176),
    to_slogic(161),
    to_slogic(169),
    to_slogic(156),
    to_slogic(156),
    to_slogic(151),
    to_slogic(151),
    to_slogic(143),
    to_slogic(116),
    to_slogic(118),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(107),
    to_slogic(119),
    to_slogic(128),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(144),
    to_slogic(118),
    to_slogic(127),
    to_slogic(134),
    to_slogic(146),
    to_slogic(141),
    to_slogic(137),
    to_slogic(134),
    to_slogic(139),
    to_slogic(151),
    to_slogic(151),
    to_slogic(149),
    to_slogic(139),
    to_slogic(110),
    to_slogic(113),
    to_slogic(121),
    to_slogic(121),
    to_slogic(101),
    to_slogic(101),
    to_slogic(103),
    to_slogic(101),
    to_slogic(134),
    to_slogic(110),
    to_slogic(143),
    to_slogic(152),
    to_slogic(157),
    to_slogic(133),
    to_slogic(110),
    to_slogic(133),
    to_slogic(133),
    to_slogic(151),
    to_slogic(155),
    to_slogic(162),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(141),
    to_slogic(151),
    to_slogic(157),
    to_slogic(155),
    to_slogic(152),
    to_slogic(133),
    to_slogic(113),
    to_slogic(87),
    to_slogic(133),
    to_slogic(157),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(176),
    to_slogic(189),
    to_slogic(177),
    to_slogic(166),
    to_slogic(185),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(193),
    to_slogic(200),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(189),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(197),
    to_slogic(204),
    to_slogic(197),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(214),
    to_slogic(205),
    to_slogic(182),
    to_slogic(166),
    to_slogic(155),
    to_slogic(130),
    to_slogic(94),
    to_slogic(82),
    to_slogic(92),
    to_slogic(101),
    to_slogic(143),
    to_slogic(191),
    to_slogic(220),
    to_slogic(171),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(64),
    to_slogic(102),
    to_slogic(141),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(151),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(96),
    to_slogic(100),
    to_slogic(92),
    to_slogic(102),
    to_slogic(99),
    to_slogic(96),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(99),
    to_slogic(115),
    to_slogic(115),
    to_slogic(135),
    to_slogic(143),
    to_slogic(156),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(152),
    to_slogic(143),
    to_slogic(121),
    to_slogic(89),
    to_slogic(81),
    to_slogic(70),
    to_slogic(76),
    to_slogic(89),
    to_slogic(89),
    to_slogic(92),
    to_slogic(100),
    to_slogic(94),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(97),
    to_slogic(100),
    to_slogic(100),
    to_slogic(97),
    to_slogic(99),
    to_slogic(89),
    to_slogic(81),
    to_slogic(99),
    to_slogic(207),
    to_slogic(205),
    to_slogic(191),
    to_slogic(197),
    to_slogic(176),
    to_slogic(172),
    to_slogic(161),
    to_slogic(156),
    to_slogic(151),
    to_slogic(151),
    to_slogic(156),
    to_slogic(143),
    to_slogic(121),
    to_slogic(116),
    to_slogic(119),
    to_slogic(124),
    to_slogic(119),
    to_slogic(128),
    to_slogic(133),
    to_slogic(125),
    to_slogic(110),
    to_slogic(119),
    to_slogic(128),
    to_slogic(137),
    to_slogic(146),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(137),
    to_slogic(110),
    to_slogic(128),
    to_slogic(133),
    to_slogic(134),
    to_slogic(139),
    to_slogic(151),
    to_slogic(128),
    to_slogic(134),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(133),
    to_slogic(110),
    to_slogic(113),
    to_slogic(133),
    to_slogic(141),
    to_slogic(133),
    to_slogic(127),
    to_slogic(117),
    to_slogic(101),
    to_slogic(96),
    to_slogic(81),
    to_slogic(96),
    to_slogic(155),
    to_slogic(162),
    to_slogic(169),
    to_slogic(155),
    to_slogic(133),
    to_slogic(122),
    to_slogic(109),
    to_slogic(118),
    to_slogic(113),
    to_slogic(110),
    to_slogic(151),
    to_slogic(152),
    to_slogic(155),
    to_slogic(143),
    to_slogic(121),
    to_slogic(121),
    to_slogic(110),
    to_slogic(134),
    to_slogic(95),
    to_slogic(119),
    to_slogic(83),
    to_slogic(63),
    to_slogic(143),
    to_slogic(157),
    to_slogic(152),
    to_slogic(182),
    to_slogic(183),
    to_slogic(166),
    to_slogic(165),
    to_slogic(182),
    to_slogic(189),
    to_slogic(193),
    to_slogic(204),
    to_slogic(200),
    to_slogic(189),
    to_slogic(193),
    to_slogic(191),
    to_slogic(196),
    to_slogic(189),
    to_slogic(196),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(197),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(204),
    to_slogic(197),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(214),
    to_slogic(213),
    to_slogic(189),
    to_slogic(156),
    to_slogic(143),
    to_slogic(102),
    to_slogic(82),
    to_slogic(82),
    to_slogic(102),
    to_slogic(102),
    to_slogic(133),
    to_slogic(182),
    to_slogic(214),
    to_slogic(213),
    to_slogic(91),
    to_slogic(33),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(50),
    to_slogic(56),
    to_slogic(81),
    to_slogic(128),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(141),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(157),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(102),
    to_slogic(96),
    to_slogic(99),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(97),
    to_slogic(109),
    to_slogic(121),
    to_slogic(135),
    to_slogic(143),
    to_slogic(151),
    to_slogic(161),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(135),
    to_slogic(121),
    to_slogic(99),
    to_slogic(76),
    to_slogic(70),
    to_slogic(81),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(97),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(97),
    to_slogic(100),
    to_slogic(97),
    to_slogic(89),
    to_slogic(76),
    to_slogic(99),
    to_slogic(207),
    to_slogic(205),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(176),
    to_slogic(169),
    to_slogic(156),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(156),
    to_slogic(130),
    to_slogic(115),
    to_slogic(116),
    to_slogic(117),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(109),
    to_slogic(119),
    to_slogic(119),
    to_slogic(146),
    to_slogic(137),
    to_slogic(139),
    to_slogic(133),
    to_slogic(137),
    to_slogic(128),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(134),
    to_slogic(139),
    to_slogic(146),
    to_slogic(149),
    to_slogic(141),
    to_slogic(128),
    to_slogic(126),
    to_slogic(149),
    to_slogic(141),
    to_slogic(117),
    to_slogic(110),
    to_slogic(102),
    to_slogic(96),
    to_slogic(81),
    to_slogic(81),
    to_slogic(69),
    to_slogic(83),
    to_slogic(143),
    to_slogic(162),
    to_slogic(162),
    to_slogic(148),
    to_slogic(127),
    to_slogic(127),
    to_slogic(126),
    to_slogic(127),
    to_slogic(102),
    to_slogic(84),
    to_slogic(84),
    to_slogic(95),
    to_slogic(89),
    to_slogic(95),
    to_slogic(81),
    to_slogic(81),
    to_slogic(71),
    to_slogic(50),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(42),
    to_slogic(110),
    to_slogic(165),
    to_slogic(182),
    to_slogic(166),
    to_slogic(162),
    to_slogic(165),
    to_slogic(185),
    to_slogic(200),
    to_slogic(189),
    to_slogic(200),
    to_slogic(200),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(189),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(197),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(213),
    to_slogic(193),
    to_slogic(177),
    to_slogic(143),
    to_slogic(118),
    to_slogic(92),
    to_slogic(75),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(125),
    to_slogic(172),
    to_slogic(196),
    to_slogic(220),
    to_slogic(143),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(63),
    to_slogic(101),
    to_slogic(141),
    to_slogic(155),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(149),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(94),
    to_slogic(94),
    to_slogic(94),
    to_slogic(102),
    to_slogic(99),
    to_slogic(100),
    to_slogic(115),
    to_slogic(115),
    to_slogic(121),
    to_slogic(135),
    to_slogic(143),
    to_slogic(156),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(161),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(100),
    to_slogic(81),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(97),
    to_slogic(97),
    to_slogic(97),
    to_slogic(89),
    to_slogic(89),
    to_slogic(82),
    to_slogic(193),
    to_slogic(205),
    to_slogic(191),
    to_slogic(197),
    to_slogic(191),
    to_slogic(183),
    to_slogic(169),
    to_slogic(143),
    to_slogic(135),
    to_slogic(121),
    to_slogic(151),
    to_slogic(143),
    to_slogic(109),
    to_slogic(102),
    to_slogic(117),
    to_slogic(119),
    to_slogic(126),
    to_slogic(117),
    to_slogic(96),
    to_slogic(119),
    to_slogic(119),
    to_slogic(139),
    to_slogic(139),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(128),
    to_slogic(119),
    to_slogic(127),
    to_slogic(125),
    to_slogic(133),
    to_slogic(133),
    to_slogic(134),
    to_slogic(127),
    to_slogic(128),
    to_slogic(141),
    to_slogic(146),
    to_slogic(134),
    to_slogic(146),
    to_slogic(117),
    to_slogic(121),
    to_slogic(141),
    to_slogic(141),
    to_slogic(117),
    to_slogic(96),
    to_slogic(101),
    to_slogic(103),
    to_slogic(87),
    to_slogic(96),
    to_slogic(88),
    to_slogic(82),
    to_slogic(103),
    to_slogic(127),
    to_slogic(141),
    to_slogic(141),
    to_slogic(136),
    to_slogic(120),
    to_slogic(89),
    to_slogic(71),
    to_slogic(76),
    to_slogic(65),
    to_slogic(91),
    to_slogic(115),
    to_slogic(71),
    to_slogic(76),
    to_slogic(58),
    to_slogic(56),
    to_slogic(50),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(42),
    to_slogic(63),
    to_slogic(148),
    to_slogic(182),
    to_slogic(162),
    to_slogic(157),
    to_slogic(177),
    to_slogic(189),
    to_slogic(200),
    to_slogic(200),
    to_slogic(193),
    to_slogic(196),
    to_slogic(193),
    to_slogic(195),
    to_slogic(196),
    to_slogic(200),
    to_slogic(193),
    to_slogic(189),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(193),
    to_slogic(162),
    to_slogic(124),
    to_slogic(107),
    to_slogic(94),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(94),
    to_slogic(96),
    to_slogic(134),
    to_slogic(158),
    to_slogic(193),
    to_slogic(213),
    to_slogic(189),
    to_slogic(64),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(75),
    to_slogic(126),
    to_slogic(151),
    to_slogic(144),
    to_slogic(141),
    to_slogic(141),
    to_slogic(149),
    to_slogic(165),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(99),
    to_slogic(94),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(94),
    to_slogic(100),
    to_slogic(109),
    to_slogic(99),
    to_slogic(109),
    to_slogic(121),
    to_slogic(135),
    to_slogic(143),
    to_slogic(156),
    to_slogic(165),
    to_slogic(169),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(144),
    to_slogic(121),
    to_slogic(92),
    to_slogic(76),
    to_slogic(70),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(89),
    to_slogic(82),
    to_slogic(176),
    to_slogic(207),
    to_slogic(205),
    to_slogic(197),
    to_slogic(197),
    to_slogic(191),
    to_slogic(169),
    to_slogic(143),
    to_slogic(121),
    to_slogic(130),
    to_slogic(135),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(128),
    to_slogic(109),
    to_slogic(110),
    to_slogic(119),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(119),
    to_slogic(133),
    to_slogic(133),
    to_slogic(134),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(146),
    to_slogic(146),
    to_slogic(134),
    to_slogic(139),
    to_slogic(117),
    to_slogic(110),
    to_slogic(141),
    to_slogic(133),
    to_slogic(121),
    to_slogic(102),
    to_slogic(121),
    to_slogic(117),
    to_slogic(110),
    to_slogic(121),
    to_slogic(133),
    to_slogic(103),
    to_slogic(82),
    to_slogic(84),
    to_slogic(97),
    to_slogic(102),
    to_slogic(126),
    to_slogic(107),
    to_slogic(82),
    to_slogic(84),
    to_slogic(65),
    to_slogic(65),
    to_slogic(97),
    to_slogic(97),
    to_slogic(71),
    to_slogic(65),
    to_slogic(71),
    to_slogic(76),
    to_slogic(49),
    to_slogic(42),
    to_slogic(36),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(102),
    to_slogic(153),
    to_slogic(177),
    to_slogic(144),
    to_slogic(155),
    to_slogic(191),
    to_slogic(204),
    to_slogic(204),
    to_slogic(193),
    to_slogic(200),
    to_slogic(189),
    to_slogic(200),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(193),
    to_slogic(196),
    to_slogic(196),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(205),
    to_slogic(204),
    to_slogic(205),
    to_slogic(205),
    to_slogic(182),
    to_slogic(143),
    to_slogic(118),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(110),
    to_slogic(125),
    to_slogic(172),
    to_slogic(189),
    to_slogic(193),
    to_slogic(193),
    to_slogic(96),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(42),
    to_slogic(50),
    to_slogic(96),
    to_slogic(139),
    to_slogic(151),
    to_slogic(151),
    to_slogic(141),
    to_slogic(151),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(121),
    to_slogic(130),
    to_slogic(143),
    to_slogic(156),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(92),
    to_slogic(81),
    to_slogic(70),
    to_slogic(81),
    to_slogic(89),
    to_slogic(92),
    to_slogic(94),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(89),
    to_slogic(97),
    to_slogic(89),
    to_slogic(77),
    to_slogic(144),
    to_slogic(213),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(191),
    to_slogic(176),
    to_slogic(143),
    to_slogic(121),
    to_slogic(109),
    to_slogic(137),
    to_slogic(139),
    to_slogic(128),
    to_slogic(117),
    to_slogic(119),
    to_slogic(119),
    to_slogic(109),
    to_slogic(101),
    to_slogic(119),
    to_slogic(128),
    to_slogic(146),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(107),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(134),
    to_slogic(133),
    to_slogic(127),
    to_slogic(119),
    to_slogic(134),
    to_slogic(146),
    to_slogic(133),
    to_slogic(134),
    to_slogic(127),
    to_slogic(117),
    to_slogic(134),
    to_slogic(133),
    to_slogic(124),
    to_slogic(113),
    to_slogic(121),
    to_slogic(128),
    to_slogic(113),
    to_slogic(102),
    to_slogic(110),
    to_slogic(88),
    to_slogic(71),
    to_slogic(63),
    to_slogic(75),
    to_slogic(69),
    to_slogic(97),
    to_slogic(107),
    to_slogic(109),
    to_slogic(91),
    to_slogic(82),
    to_slogic(91),
    to_slogic(102),
    to_slogic(83),
    to_slogic(84),
    to_slogic(76),
    to_slogic(58),
    to_slogic(81),
    to_slogic(71),
    to_slogic(50),
    to_slogic(40),
    to_slogic(36),
    to_slogic(36),
    to_slogic(42),
    to_slogic(102),
    to_slogic(170),
    to_slogic(158),
    to_slogic(139),
    to_slogic(162),
    to_slogic(182),
    to_slogic(200),
    to_slogic(193),
    to_slogic(200),
    to_slogic(196),
    to_slogic(196),
    to_slogic(189),
    to_slogic(196),
    to_slogic(193),
    to_slogic(189),
    to_slogic(196),
    to_slogic(196),
    to_slogic(189),
    to_slogic(196),
    to_slogic(193),
    to_slogic(196),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(196),
    to_slogic(204),
    to_slogic(205),
    to_slogic(204),
    to_slogic(189),
    to_slogic(136),
    to_slogic(96),
    to_slogic(88),
    to_slogic(82),
    to_slogic(89),
    to_slogic(82),
    to_slogic(94),
    to_slogic(94),
    to_slogic(96),
    to_slogic(101),
    to_slogic(119),
    to_slogic(149),
    to_slogic(172),
    to_slogic(193),
    to_slogic(198),
    to_slogic(144),
    to_slogic(64),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(40),
    to_slogic(42),
    to_slogic(63),
    to_slogic(121),
    to_slogic(151),
    to_slogic(143),
    to_slogic(141),
    to_slogic(151),
    to_slogic(149),
    to_slogic(165),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(150),
    to_slogic(100),
    to_slogic(101),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(99),
    to_slogic(115),
    to_slogic(121),
    to_slogic(135),
    to_slogic(143),
    to_slogic(157),
    to_slogic(161),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(143),
    to_slogic(121),
    to_slogic(99),
    to_slogic(75),
    to_slogic(76),
    to_slogic(81),
    to_slogic(81),
    to_slogic(92),
    to_slogic(97),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(97),
    to_slogic(100),
    to_slogic(100),
    to_slogic(97),
    to_slogic(99),
    to_slogic(97),
    to_slogic(89),
    to_slogic(89),
    to_slogic(81),
    to_slogic(121),
    to_slogic(213),
    to_slogic(203),
    to_slogic(205),
    to_slogic(197),
    to_slogic(197),
    to_slogic(172),
    to_slogic(143),
    to_slogic(121),
    to_slogic(126),
    to_slogic(157),
    to_slogic(137),
    to_slogic(144),
    to_slogic(117),
    to_slogic(119),
    to_slogic(109),
    to_slogic(102),
    to_slogic(119),
    to_slogic(128),
    to_slogic(139),
    to_slogic(133),
    to_slogic(146),
    to_slogic(133),
    to_slogic(127),
    to_slogic(119),
    to_slogic(127),
    to_slogic(128),
    to_slogic(133),
    to_slogic(134),
    to_slogic(133),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(117),
    to_slogic(101),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(110),
    to_slogic(113),
    to_slogic(122),
    to_slogic(102),
    to_slogic(96),
    to_slogic(75),
    to_slogic(63),
    to_slogic(50),
    to_slogic(64),
    to_slogic(50),
    to_slogic(64),
    to_slogic(82),
    to_slogic(103),
    to_slogic(117),
    to_slogic(102),
    to_slogic(102),
    to_slogic(89),
    to_slogic(118),
    to_slogic(84),
    to_slogic(120),
    to_slogic(71),
    to_slogic(65),
    to_slogic(58),
    to_slogic(81),
    to_slogic(84),
    to_slogic(42),
    to_slogic(42),
    to_slogic(42),
    to_slogic(58),
    to_slogic(119),
    to_slogic(176),
    to_slogic(143),
    to_slogic(127),
    to_slogic(158),
    to_slogic(193),
    to_slogic(189),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(196),
    to_slogic(193),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(167),
    to_slogic(109),
    to_slogic(92),
    to_slogic(94),
    to_slogic(92),
    to_slogic(96),
    to_slogic(82),
    to_slogic(92),
    to_slogic(96),
    to_slogic(110),
    to_slogic(120),
    to_slogic(141),
    to_slogic(162),
    to_slogic(182),
    to_slogic(198),
    to_slogic(193),
    to_slogic(149),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(50),
    to_slogic(56),
    to_slogic(87),
    to_slogic(132),
    to_slogic(151),
    to_slogic(144),
    to_slogic(141),
    to_slogic(151),
    to_slogic(155),
    to_slogic(166),
    to_slogic(165),
    to_slogic(162),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(115),
    to_slogic(109),
    to_slogic(121),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(161),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(99),
    to_slogic(81),
    to_slogic(70),
    to_slogic(81),
    to_slogic(82),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(89),
    to_slogic(100),
    to_slogic(100),
    to_slogic(97),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(97),
    to_slogic(100),
    to_slogic(97),
    to_slogic(100),
    to_slogic(81),
    to_slogic(92),
    to_slogic(207),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(196),
    to_slogic(176),
    to_slogic(143),
    to_slogic(130),
    to_slogic(144),
    to_slogic(137),
    to_slogic(146),
    to_slogic(133),
    to_slogic(133),
    to_slogic(109),
    to_slogic(101),
    to_slogic(110),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(134),
    to_slogic(133),
    to_slogic(127),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(133),
    to_slogic(127),
    to_slogic(119),
    to_slogic(134),
    to_slogic(146),
    to_slogic(133),
    to_slogic(134),
    to_slogic(124),
    to_slogic(101),
    to_slogic(133),
    to_slogic(127),
    to_slogic(134),
    to_slogic(128),
    to_slogic(96),
    to_slogic(88),
    to_slogic(71),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(69),
    to_slogic(50),
    to_slogic(64),
    to_slogic(50),
    to_slogic(76),
    to_slogic(109),
    to_slogic(102),
    to_slogic(107),
    to_slogic(84),
    to_slogic(63),
    to_slogic(65),
    to_slogic(89),
    to_slogic(97),
    to_slogic(89),
    to_slogic(84),
    to_slogic(78),
    to_slogic(50),
    to_slogic(81),
    to_slogic(76),
    to_slogic(36),
    to_slogic(36),
    to_slogic(63),
    to_slogic(133),
    to_slogic(170),
    to_slogic(137),
    to_slogic(120),
    to_slogic(158),
    to_slogic(189),
    to_slogic(198),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(182),
    to_slogic(196),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(191),
    to_slogic(193),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(193),
    to_slogic(158),
    to_slogic(119),
    to_slogic(133),
    to_slogic(120),
    to_slogic(96),
    to_slogic(96),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(110),
    to_slogic(139),
    to_slogic(152),
    to_slogic(162),
    to_slogic(162),
    to_slogic(177),
    to_slogic(183),
    to_slogic(193),
    to_slogic(166),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(120),
    to_slogic(141),
    to_slogic(151),
    to_slogic(151),
    to_slogic(143),
    to_slogic(162),
    to_slogic(165),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(158),
    to_slogic(162),
    to_slogic(156),
    to_slogic(149),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(149),
    to_slogic(155),
    to_slogic(150),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(97),
    to_slogic(109),
    to_slogic(121),
    to_slogic(135),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(94),
    to_slogic(82),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(97),
    to_slogic(99),
    to_slogic(100),
    to_slogic(89),
    to_slogic(81),
    to_slogic(76),
    to_slogic(178),
    to_slogic(207),
    to_slogic(205),
    to_slogic(183),
    to_slogic(197),
    to_slogic(176),
    to_slogic(161),
    to_slogic(130),
    to_slogic(118),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(119),
    to_slogic(102),
    to_slogic(110),
    to_slogic(119),
    to_slogic(133),
    to_slogic(134),
    to_slogic(133),
    to_slogic(139),
    to_slogic(119),
    to_slogic(119),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(128),
    to_slogic(119),
    to_slogic(128),
    to_slogic(146),
    to_slogic(146),
    to_slogic(133),
    to_slogic(128),
    to_slogic(127),
    to_slogic(103),
    to_slogic(141),
    to_slogic(127),
    to_slogic(110),
    to_slogic(82),
    to_slogic(69),
    to_slogic(69),
    to_slogic(88),
    to_slogic(91),
    to_slogic(75),
    to_slogic(64),
    to_slogic(56),
    to_slogic(46),
    to_slogic(50),
    to_slogic(50),
    to_slogic(103),
    to_slogic(122),
    to_slogic(115),
    to_slogic(88),
    to_slogic(46),
    to_slogic(46),
    to_slogic(71),
    to_slogic(107),
    to_slogic(65),
    to_slogic(97),
    to_slogic(89),
    to_slogic(50),
    to_slogic(42),
    to_slogic(89),
    to_slogic(71),
    to_slogic(40),
    to_slogic(63),
    to_slogic(143),
    to_slogic(166),
    to_slogic(133),
    to_slogic(141),
    to_slogic(170),
    to_slogic(193),
    to_slogic(198),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(185),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(182),
    to_slogic(189),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(196),
    to_slogic(171),
    to_slogic(109),
    to_slogic(102),
    to_slogic(110),
    to_slogic(134),
    to_slogic(133),
    to_slogic(119),
    to_slogic(101),
    to_slogic(110),
    to_slogic(128),
    to_slogic(151),
    to_slogic(157),
    to_slogic(162),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(177),
    to_slogic(193),
    to_slogic(166),
    to_slogic(64),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(87),
    to_slogic(133),
    to_slogic(151),
    to_slogic(151),
    to_slogic(139),
    to_slogic(151),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(158),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(162),
    to_slogic(156),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(151),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(96),
    to_slogic(100),
    to_slogic(109),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(115),
    to_slogic(121),
    to_slogic(130),
    to_slogic(143),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(156),
    to_slogic(143),
    to_slogic(121),
    to_slogic(100),
    to_slogic(81),
    to_slogic(70),
    to_slogic(76),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(97),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(76),
    to_slogic(126),
    to_slogic(213),
    to_slogic(197),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(165),
    to_slogic(157),
    to_slogic(137),
    to_slogic(144),
    to_slogic(137),
    to_slogic(130),
    to_slogic(117),
    to_slogic(109),
    to_slogic(124),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(119),
    to_slogic(110),
    to_slogic(119),
    to_slogic(128),
    to_slogic(134),
    to_slogic(128),
    to_slogic(119),
    to_slogic(128),
    to_slogic(119),
    to_slogic(117),
    to_slogic(146),
    to_slogic(127),
    to_slogic(133),
    to_slogic(134),
    to_slogic(149),
    to_slogic(126),
    to_slogic(103),
    to_slogic(133),
    to_slogic(96),
    to_slogic(75),
    to_slogic(56),
    to_slogic(69),
    to_slogic(91),
    to_slogic(81),
    to_slogic(56),
    to_slogic(46),
    to_slogic(50),
    to_slogic(49),
    to_slogic(50),
    to_slogic(50),
    to_slogic(82),
    to_slogic(122),
    to_slogic(113),
    to_slogic(81),
    to_slogic(50),
    to_slogic(50),
    to_slogic(69),
    to_slogic(115),
    to_slogic(76),
    to_slogic(84),
    to_slogic(89),
    to_slogic(50),
    to_slogic(42),
    to_slogic(42),
    to_slogic(102),
    to_slogic(84),
    to_slogic(71),
    to_slogic(149),
    to_slogic(162),
    to_slogic(125),
    to_slogic(141),
    to_slogic(185),
    to_slogic(200),
    to_slogic(189),
    to_slogic(182),
    to_slogic(182),
    to_slogic(177),
    to_slogic(182),
    to_slogic(189),
    to_slogic(185),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(182),
    to_slogic(185),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(196),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(193),
    to_slogic(171),
    to_slogic(118),
    to_slogic(96),
    to_slogic(81),
    to_slogic(102),
    to_slogic(102),
    to_slogic(134),
    to_slogic(141),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(173),
    to_slogic(165),
    to_slogic(177),
    to_slogic(198),
    to_slogic(166),
    to_slogic(62),
    to_slogic(33),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(64),
    to_slogic(110),
    to_slogic(141),
    to_slogic(143),
    to_slogic(151),
    to_slogic(141),
    to_slogic(149),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(167),
    to_slogic(162),
    to_slogic(167),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(158),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(149),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(99),
    to_slogic(109),
    to_slogic(121),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(161),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(92),
    to_slogic(81),
    to_slogic(70),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(97),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(82),
    to_slogic(109),
    to_slogic(207),
    to_slogic(205),
    to_slogic(191),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(157),
    to_slogic(165),
    to_slogic(144),
    to_slogic(157),
    to_slogic(115),
    to_slogic(101),
    to_slogic(119),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(134),
    to_slogic(119),
    to_slogic(102),
    to_slogic(119),
    to_slogic(126),
    to_slogic(127),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(119),
    to_slogic(119),
    to_slogic(133),
    to_slogic(120),
    to_slogic(101),
    to_slogic(110),
    to_slogic(128),
    to_slogic(149),
    to_slogic(134),
    to_slogic(103),
    to_slogic(96),
    to_slogic(63),
    to_slogic(63),
    to_slogic(75),
    to_slogic(84),
    to_slogic(63),
    to_slogic(50),
    to_slogic(46),
    to_slogic(56),
    to_slogic(56),
    to_slogic(46),
    to_slogic(46),
    to_slogic(50),
    to_slogic(107),
    to_slogic(102),
    to_slogic(81),
    to_slogic(50),
    to_slogic(46),
    to_slogic(76),
    to_slogic(115),
    to_slogic(102),
    to_slogic(84),
    to_slogic(97),
    to_slogic(42),
    to_slogic(50),
    to_slogic(58),
    to_slogic(42),
    to_slogic(102),
    to_slogic(95),
    to_slogic(149),
    to_slogic(158),
    to_slogic(128),
    to_slogic(144),
    to_slogic(176),
    to_slogic(193),
    to_slogic(193),
    to_slogic(182),
    to_slogic(185),
    to_slogic(176),
    to_slogic(182),
    to_slogic(185),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(185),
    to_slogic(185),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(204),
    to_slogic(193),
    to_slogic(176),
    to_slogic(124),
    to_slogic(83),
    to_slogic(56),
    to_slogic(102),
    to_slogic(110),
    to_slogic(102),
    to_slogic(110),
    to_slogic(126),
    to_slogic(143),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(162),
    to_slogic(173),
    to_slogic(172),
    to_slogic(183),
    to_slogic(207),
    to_slogic(171),
    to_slogic(75),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(75),
    to_slogic(125),
    to_slogic(151),
    to_slogic(151),
    to_slogic(139),
    to_slogic(151),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(162),
    to_slogic(166),
    to_slogic(165),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(149),
    to_slogic(155),
    to_slogic(156),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(97),
    to_slogic(109),
    to_slogic(121),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(143),
    to_slogic(130),
    to_slogic(100),
    to_slogic(81),
    to_slogic(76),
    to_slogic(75),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(94),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(89),
    to_slogic(178),
    to_slogic(207),
    to_slogic(205),
    to_slogic(191),
    to_slogic(191),
    to_slogic(165),
    to_slogic(178),
    to_slogic(173),
    to_slogic(157),
    to_slogic(143),
    to_slogic(109),
    to_slogic(109),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(133),
    to_slogic(128),
    to_slogic(117),
    to_slogic(109),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(119),
    to_slogic(128),
    to_slogic(127),
    to_slogic(117),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(128),
    to_slogic(110),
    to_slogic(87),
    to_slogic(103),
    to_slogic(119),
    to_slogic(81),
    to_slogic(63),
    to_slogic(65),
    to_slogic(83),
    to_slogic(75),
    to_slogic(69),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(69),
    to_slogic(44),
    to_slogic(40),
    to_slogic(46),
    to_slogic(84),
    to_slogic(102),
    to_slogic(64),
    to_slogic(56),
    to_slogic(50),
    to_slogic(63),
    to_slogic(102),
    to_slogic(84),
    to_slogic(103),
    to_slogic(115),
    to_slogic(63),
    to_slogic(50),
    to_slogic(109),
    to_slogic(44),
    to_slogic(56),
    to_slogic(130),
    to_slogic(158),
    to_slogic(137),
    to_slogic(127),
    to_slogic(144),
    to_slogic(189),
    to_slogic(193),
    to_slogic(200),
    to_slogic(189),
    to_slogic(185),
    to_slogic(176),
    to_slogic(182),
    to_slogic(177),
    to_slogic(185),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(170),
    to_slogic(182),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(193),
    to_slogic(196),
    to_slogic(189),
    to_slogic(166),
    to_slogic(82),
    to_slogic(56),
    to_slogic(101),
    to_slogic(81),
    to_slogic(101),
    to_slogic(134),
    to_slogic(110),
    to_slogic(121),
    to_slogic(110),
    to_slogic(143),
    to_slogic(157),
    to_slogic(155),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(187),
    to_slogic(198),
    to_slogic(183),
    to_slogic(64),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(64),
    to_slogic(96),
    to_slogic(139),
    to_slogic(151),
    to_slogic(139),
    to_slogic(141),
    to_slogic(155),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(166),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(157),
    to_slogic(162),
    to_slogic(157),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(109),
    to_slogic(109),
    to_slogic(96),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(97),
    to_slogic(115),
    to_slogic(130),
    to_slogic(143),
    to_slogic(156),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(152),
    to_slogic(144),
    to_slogic(121),
    to_slogic(100),
    to_slogic(76),
    to_slogic(63),
    to_slogic(81),
    to_slogic(82),
    to_slogic(89),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(89),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(82),
    to_slogic(121),
    to_slogic(207),
    to_slogic(207),
    to_slogic(205),
    to_slogic(191),
    to_slogic(165),
    to_slogic(165),
    to_slogic(178),
    to_slogic(158),
    to_slogic(117),
    to_slogic(92),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(109),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(119),
    to_slogic(119),
    to_slogic(119),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(146),
    to_slogic(134),
    to_slogic(117),
    to_slogic(82),
    to_slogic(83),
    to_slogic(81),
    to_slogic(75),
    to_slogic(83),
    to_slogic(75),
    to_slogic(82),
    to_slogic(84),
    to_slogic(71),
    to_slogic(65),
    to_slogic(50),
    to_slogic(50),
    to_slogic(97),
    to_slogic(64),
    to_slogic(42),
    to_slogic(36),
    to_slogic(65),
    to_slogic(81),
    to_slogic(89),
    to_slogic(46),
    to_slogic(46),
    to_slogic(50),
    to_slogic(81),
    to_slogic(84),
    to_slogic(82),
    to_slogic(97),
    to_slogic(71),
    to_slogic(44),
    to_slogic(109),
    to_slogic(97),
    to_slogic(36),
    to_slogic(107),
    to_slogic(162),
    to_slogic(139),
    to_slogic(120),
    to_slogic(144),
    to_slogic(189),
    to_slogic(200),
    to_slogic(193),
    to_slogic(189),
    to_slogic(189),
    to_slogic(185),
    to_slogic(182),
    to_slogic(177),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(182),
    to_slogic(170),
    to_slogic(176),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(185),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(189),
    to_slogic(193),
    to_slogic(189),
    to_slogic(155),
    to_slogic(82),
    to_slogic(64),
    to_slogic(56),
    to_slogic(91),
    to_slogic(102),
    to_slogic(81),
    to_slogic(126),
    to_slogic(126),
    to_slogic(119),
    to_slogic(113),
    to_slogic(133),
    to_slogic(152),
    to_slogic(155),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(183),
    to_slogic(198),
    to_slogic(136),
    to_slogic(62),
    to_slogic(40),
    to_slogic(33),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(68),
    to_slogic(117),
    to_slogic(139),
    to_slogic(141),
    to_slogic(139),
    to_slogic(151),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(166),
    to_slogic(165),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(162),
    to_slogic(155),
    to_slogic(158),
    to_slogic(149),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(100),
    to_slogic(99),
    to_slogic(94),
    to_slogic(100),
    to_slogic(97),
    to_slogic(121),
    to_slogic(121),
    to_slogic(143),
    to_slogic(152),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(157),
    to_slogic(156),
    to_slogic(143),
    to_slogic(121),
    to_slogic(99),
    to_slogic(81),
    to_slogic(70),
    to_slogic(76),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(97),
    to_slogic(92),
    to_slogic(97),
    to_slogic(99),
    to_slogic(97),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(89),
    to_slogic(158),
    to_slogic(213),
    to_slogic(207),
    to_slogic(197),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(116),
    to_slogic(117),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(128),
    to_slogic(117),
    to_slogic(110),
    to_slogic(128),
    to_slogic(128),
    to_slogic(127),
    to_slogic(128),
    to_slogic(119),
    to_slogic(124),
    to_slogic(119),
    to_slogic(124),
    to_slogic(134),
    to_slogic(128),
    to_slogic(119),
    to_slogic(110),
    to_slogic(101),
    to_slogic(88),
    to_slogic(69),
    to_slogic(69),
    to_slogic(75),
    to_slogic(65),
    to_slogic(83),
    to_slogic(81),
    to_slogic(69),
    to_slogic(56),
    to_slogic(50),
    to_slogic(46),
    to_slogic(83),
    to_slogic(102),
    to_slogic(40),
    to_slogic(36),
    to_slogic(46),
    to_slogic(82),
    to_slogic(75),
    to_slogic(69),
    to_slogic(44),
    to_slogic(50),
    to_slogic(64),
    to_slogic(63),
    to_slogic(50),
    to_slogic(56),
    to_slogic(97),
    to_slogic(44),
    to_slogic(58),
    to_slogic(145),
    to_slogic(65),
    to_slogic(71),
    to_slogic(127),
    to_slogic(117),
    to_slogic(121),
    to_slogic(158),
    to_slogic(195),
    to_slogic(193),
    to_slogic(200),
    to_slogic(189),
    to_slogic(189),
    to_slogic(189),
    to_slogic(176),
    to_slogic(185),
    to_slogic(182),
    to_slogic(177),
    to_slogic(185),
    to_slogic(182),
    to_slogic(170),
    to_slogic(171),
    to_slogic(176),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(189),
    to_slogic(185),
    to_slogic(193),
    to_slogic(176),
    to_slogic(155),
    to_slogic(102),
    to_slogic(75),
    to_slogic(96),
    to_slogic(75),
    to_slogic(101),
    to_slogic(101),
    to_slogic(89),
    to_slogic(133),
    to_slogic(121),
    to_slogic(121),
    to_slogic(110),
    to_slogic(149),
    to_slogic(151),
    to_slogic(162),
    to_slogic(173),
    to_slogic(178),
    to_slogic(193),
    to_slogic(191),
    to_slogic(102),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(87),
    to_slogic(125),
    to_slogic(133),
    to_slogic(139),
    to_slogic(134),
    to_slogic(144),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(156),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(97),
    to_slogic(100),
    to_slogic(115),
    to_slogic(130),
    to_slogic(143),
    to_slogic(156),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(143),
    to_slogic(130),
    to_slogic(92),
    to_slogic(76),
    to_slogic(70),
    to_slogic(82),
    to_slogic(82),
    to_slogic(89),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(100),
    to_slogic(191),
    to_slogic(213),
    to_slogic(197),
    to_slogic(191),
    to_slogic(183),
    to_slogic(183),
    to_slogic(165),
    to_slogic(116),
    to_slogic(137),
    to_slogic(124),
    to_slogic(128),
    to_slogic(127),
    to_slogic(119),
    to_slogic(117),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(127),
    to_slogic(121),
    to_slogic(121),
    to_slogic(117),
    to_slogic(133),
    to_slogic(128),
    to_slogic(124),
    to_slogic(117),
    to_slogic(117),
    to_slogic(110),
    to_slogic(103),
    to_slogic(103),
    to_slogic(81),
    to_slogic(65),
    to_slogic(82),
    to_slogic(89),
    to_slogic(65),
    to_slogic(50),
    to_slogic(42),
    to_slogic(36),
    to_slogic(63),
    to_slogic(102),
    to_slogic(97),
    to_slogic(44),
    to_slogic(46),
    to_slogic(46),
    to_slogic(75),
    to_slogic(75),
    to_slogic(69),
    to_slogic(46),
    to_slogic(64),
    to_slogic(46),
    to_slogic(50),
    to_slogic(50),
    to_slogic(63),
    to_slogic(103),
    to_slogic(42),
    to_slogic(84),
    to_slogic(122),
    to_slogic(102),
    to_slogic(127),
    to_slogic(102),
    to_slogic(101),
    to_slogic(148),
    to_slogic(189),
    to_slogic(193),
    to_slogic(193),
    to_slogic(189),
    to_slogic(191),
    to_slogic(185),
    to_slogic(185),
    to_slogic(185),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(176),
    to_slogic(165),
    to_slogic(176),
    to_slogic(185),
    to_slogic(176),
    to_slogic(185),
    to_slogic(185),
    to_slogic(189),
    to_slogic(185),
    to_slogic(179),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(172),
    to_slogic(127),
    to_slogic(92),
    to_slogic(77),
    to_slogic(102),
    to_slogic(96),
    to_slogic(95),
    to_slogic(102),
    to_slogic(114),
    to_slogic(127),
    to_slogic(126),
    to_slogic(107),
    to_slogic(141),
    to_slogic(157),
    to_slogic(173),
    to_slogic(183),
    to_slogic(193),
    to_slogic(172),
    to_slogic(94),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(69),
    to_slogic(101),
    to_slogic(132),
    to_slogic(134),
    to_slogic(125),
    to_slogic(134),
    to_slogic(156),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(156),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(149),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(97),
    to_slogic(109),
    to_slogic(130),
    to_slogic(135),
    to_slogic(152),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(99),
    to_slogic(81),
    to_slogic(76),
    to_slogic(75),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(99),
    to_slogic(82),
    to_slogic(144),
    to_slogic(213),
    to_slogic(197),
    to_slogic(191),
    to_slogic(183),
    to_slogic(197),
    to_slogic(133),
    to_slogic(126),
    to_slogic(144),
    to_slogic(109),
    to_slogic(124),
    to_slogic(128),
    to_slogic(119),
    to_slogic(119),
    to_slogic(128),
    to_slogic(127),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(121),
    to_slogic(133),
    to_slogic(122),
    to_slogic(113),
    to_slogic(113),
    to_slogic(128),
    to_slogic(121),
    to_slogic(103),
    to_slogic(69),
    to_slogic(81),
    to_slogic(69),
    to_slogic(81),
    to_slogic(82),
    to_slogic(96),
    to_slogic(96),
    to_slogic(56),
    to_slogic(50),
    to_slogic(49),
    to_slogic(42),
    to_slogic(63),
    to_slogic(107),
    to_slogic(75),
    to_slogic(36),
    to_slogic(49),
    to_slogic(75),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(75),
    to_slogic(76),
    to_slogic(76),
    to_slogic(63),
    to_slogic(76),
    to_slogic(91),
    to_slogic(63),
    to_slogic(109),
    to_slogic(107),
    to_slogic(133),
    to_slogic(136),
    to_slogic(102),
    to_slogic(148),
    to_slogic(166),
    to_slogic(193),
    to_slogic(189),
    to_slogic(185),
    to_slogic(193),
    to_slogic(189),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(170),
    to_slogic(176),
    to_slogic(170),
    to_slogic(185),
    to_slogic(185),
    to_slogic(185),
    to_slogic(185),
    to_slogic(185),
    to_slogic(185),
    to_slogic(185),
    to_slogic(187),
    to_slogic(195),
    to_slogic(193),
    to_slogic(195),
    to_slogic(187),
    to_slogic(151),
    to_slogic(115),
    to_slogic(81),
    to_slogic(82),
    to_slogic(121),
    to_slogic(110),
    to_slogic(101),
    to_slogic(96),
    to_slogic(133),
    to_slogic(133),
    to_slogic(126),
    to_slogic(141),
    to_slogic(157),
    to_slogic(182),
    to_slogic(183),
    to_slogic(130),
    to_slogic(64),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(83),
    to_slogic(120),
    to_slogic(132),
    to_slogic(125),
    to_slogic(125),
    to_slogic(141),
    to_slogic(156),
    to_slogic(172),
    to_slogic(166),
    to_slogic(172),
    to_slogic(166),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(166),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(158),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(99),
    to_slogic(99),
    to_slogic(97),
    to_slogic(109),
    to_slogic(121),
    to_slogic(143),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(143),
    to_slogic(130),
    to_slogic(99),
    to_slogic(76),
    to_slogic(62),
    to_slogic(76),
    to_slogic(81),
    to_slogic(89),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(97),
    to_slogic(99),
    to_slogic(94),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(102),
    to_slogic(198),
    to_slogic(207),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(144),
    to_slogic(143),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(110),
    to_slogic(101),
    to_slogic(127),
    to_slogic(128),
    to_slogic(127),
    to_slogic(119),
    to_slogic(119),
    to_slogic(110),
    to_slogic(126),
    to_slogic(127),
    to_slogic(128),
    to_slogic(127),
    to_slogic(133),
    to_slogic(113),
    to_slogic(88),
    to_slogic(69),
    to_slogic(69),
    to_slogic(69),
    to_slogic(75),
    to_slogic(81),
    to_slogic(88),
    to_slogic(91),
    to_slogic(75),
    to_slogic(63),
    to_slogic(56),
    to_slogic(50),
    to_slogic(46),
    to_slogic(65),
    to_slogic(88),
    to_slogic(81),
    to_slogic(50),
    to_slogic(63),
    to_slogic(75),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(68),
    to_slogic(65),
    to_slogic(56),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(91),
    to_slogic(91),
    to_slogic(115),
    to_slogic(126),
    to_slogic(143),
    to_slogic(171),
    to_slogic(177),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(185),
    to_slogic(185),
    to_slogic(182),
    to_slogic(170),
    to_slogic(176),
    to_slogic(182),
    to_slogic(170),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(182),
    to_slogic(170),
    to_slogic(176),
    to_slogic(177),
    to_slogic(185),
    to_slogic(185),
    to_slogic(193),
    to_slogic(195),
    to_slogic(187),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(193),
    to_slogic(165),
    to_slogic(134),
    to_slogic(99),
    to_slogic(83),
    to_slogic(69),
    to_slogic(102),
    to_slogic(89),
    to_slogic(81),
    to_slogic(95),
    to_slogic(134),
    to_slogic(134),
    to_slogic(133),
    to_slogic(157),
    to_slogic(157),
    to_slogic(118),
    to_slogic(70),
    to_slogic(44),
    to_slogic(36),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(69),
    to_slogic(96),
    to_slogic(125),
    to_slogic(132),
    to_slogic(125),
    to_slogic(134),
    to_slogic(144),
    to_slogic(172),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(156),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(166),
    to_slogic(165),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(94),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(92),
    to_slogic(89),
    to_slogic(100),
    to_slogic(130),
    to_slogic(143),
    to_slogic(151),
    to_slogic(157),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(152),
    to_slogic(143),
    to_slogic(130),
    to_slogic(100),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(183),
    to_slogic(222),
    to_slogic(205),
    to_slogic(197),
    to_slogic(197),
    to_slogic(165),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(119),
    to_slogic(102),
    to_slogic(110),
    to_slogic(127),
    to_slogic(128),
    to_slogic(119),
    to_slogic(117),
    to_slogic(110),
    to_slogic(133),
    to_slogic(127),
    to_slogic(127),
    to_slogic(124),
    to_slogic(103),
    to_slogic(133),
    to_slogic(127),
    to_slogic(87),
    to_slogic(69),
    to_slogic(71),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(81),
    to_slogic(89),
    to_slogic(75),
    to_slogic(63),
    to_slogic(50),
    to_slogic(50),
    to_slogic(56),
    to_slogic(69),
    to_slogic(63),
    to_slogic(91),
    to_slogic(84),
    to_slogic(63),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(75),
    to_slogic(89),
    to_slogic(84),
    to_slogic(78),
    to_slogic(109),
    to_slogic(120),
    to_slogic(143),
    to_slogic(153),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(177),
    to_slogic(182),
    to_slogic(176),
    to_slogic(170),
    to_slogic(167),
    to_slogic(165),
    to_slogic(176),
    to_slogic(170),
    to_slogic(176),
    to_slogic(170),
    to_slogic(176),
    to_slogic(170),
    to_slogic(170),
    to_slogic(176),
    to_slogic(176),
    to_slogic(185),
    to_slogic(195),
    to_slogic(193),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(193),
    to_slogic(187),
    to_slogic(146),
    to_slogic(115),
    to_slogic(82),
    to_slogic(69),
    to_slogic(64),
    to_slogic(102),
    to_slogic(87),
    to_slogic(69),
    to_slogic(126),
    to_slogic(134),
    to_slogic(142),
    to_slogic(149),
    to_slogic(139),
    to_slogic(116),
    to_slogic(63),
    to_slogic(44),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(75),
    to_slogic(120),
    to_slogic(139),
    to_slogic(125),
    to_slogic(127),
    to_slogic(130),
    to_slogic(149),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(156),
    to_slogic(165),
    to_slogic(166),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(92),
    to_slogic(109),
    to_slogic(121),
    to_slogic(143),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(143),
    to_slogic(121),
    to_slogic(100),
    to_slogic(76),
    to_slogic(63),
    to_slogic(81),
    to_slogic(77),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(99),
    to_slogic(102),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(92),
    to_slogic(92),
    to_slogic(187),
    to_slogic(213),
    to_slogic(213),
    to_slogic(205),
    to_slogic(191),
    to_slogic(151),
    to_slogic(116),
    to_slogic(126),
    to_slogic(119),
    to_slogic(119),
    to_slogic(110),
    to_slogic(128),
    to_slogic(128),
    to_slogic(110),
    to_slogic(117),
    to_slogic(128),
    to_slogic(134),
    to_slogic(134),
    to_slogic(128),
    to_slogic(128),
    to_slogic(110),
    to_slogic(96),
    to_slogic(110),
    to_slogic(81),
    to_slogic(81),
    to_slogic(75),
    to_slogic(63),
    to_slogic(56),
    to_slogic(50),
    to_slogic(50),
    to_slogic(69),
    to_slogic(75),
    to_slogic(69),
    to_slogic(71),
    to_slogic(75),
    to_slogic(63),
    to_slogic(50),
    to_slogic(76),
    to_slogic(50),
    to_slogic(102),
    to_slogic(107),
    to_slogic(69),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(42),
    to_slogic(63),
    to_slogic(102),
    to_slogic(103),
    to_slogic(88),
    to_slogic(91),
    to_slogic(145),
    to_slogic(148),
    to_slogic(170),
    to_slogic(167),
    to_slogic(176),
    to_slogic(176),
    to_slogic(185),
    to_slogic(189),
    to_slogic(182),
    to_slogic(170),
    to_slogic(167),
    to_slogic(172),
    to_slogic(170),
    to_slogic(177),
    to_slogic(176),
    to_slogic(176),
    to_slogic(172),
    to_slogic(170),
    to_slogic(176),
    to_slogic(172),
    to_slogic(176),
    to_slogic(193),
    to_slogic(193),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(187),
    to_slogic(157),
    to_slogic(118),
    to_slogic(89),
    to_slogic(77),
    to_slogic(49),
    to_slogic(49),
    to_slogic(101),
    to_slogic(75),
    to_slogic(96),
    to_slogic(134),
    to_slogic(134),
    to_slogic(157),
    to_slogic(141),
    to_slogic(116),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(33),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(64),
    to_slogic(96),
    to_slogic(125),
    to_slogic(132),
    to_slogic(125),
    to_slogic(120),
    to_slogic(141),
    to_slogic(156),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(166),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(166),
    to_slogic(162),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(97),
    to_slogic(92),
    to_slogic(109),
    to_slogic(124),
    to_slogic(135),
    to_slogic(152),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(144),
    to_slogic(130),
    to_slogic(100),
    to_slogic(76),
    to_slogic(70),
    to_slogic(77),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(92),
    to_slogic(99),
    to_slogic(187),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(175),
    to_slogic(115),
    to_slogic(109),
    to_slogic(128),
    to_slogic(119),
    to_slogic(119),
    to_slogic(126),
    to_slogic(119),
    to_slogic(110),
    to_slogic(109),
    to_slogic(128),
    to_slogic(127),
    to_slogic(139),
    to_slogic(134),
    to_slogic(128),
    to_slogic(124),
    to_slogic(101),
    to_slogic(77),
    to_slogic(76),
    to_slogic(56),
    to_slogic(75),
    to_slogic(81),
    to_slogic(50),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(84),
    to_slogic(69),
    to_slogic(71),
    to_slogic(88),
    to_slogic(56),
    to_slogic(50),
    to_slogic(71),
    to_slogic(46),
    to_slogic(78),
    to_slogic(127),
    to_slogic(91),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(36),
    to_slogic(50),
    to_slogic(101),
    to_slogic(113),
    to_slogic(83),
    to_slogic(113),
    to_slogic(127),
    to_slogic(160),
    to_slogic(162),
    to_slogic(182),
    to_slogic(182),
    to_slogic(182),
    to_slogic(185),
    to_slogic(189),
    to_slogic(182),
    to_slogic(170),
    to_slogic(167),
    to_slogic(158),
    to_slogic(165),
    to_slogic(172),
    to_slogic(176),
    to_slogic(176),
    to_slogic(176),
    to_slogic(156),
    to_slogic(162),
    to_slogic(172),
    to_slogic(176),
    to_slogic(187),
    to_slogic(195),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(195),
    to_slogic(195),
    to_slogic(195),
    to_slogic(200),
    to_slogic(195),
    to_slogic(200),
    to_slogic(193),
    to_slogic(179),
    to_slogic(165),
    to_slogic(126),
    to_slogic(97),
    to_slogic(76),
    to_slogic(49),
    to_slogic(44),
    to_slogic(75),
    to_slogic(81),
    to_slogic(81),
    to_slogic(133),
    to_slogic(134),
    to_slogic(157),
    to_slogic(141),
    to_slogic(102),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(68),
    to_slogic(109),
    to_slogic(141),
    to_slogic(130),
    to_slogic(125),
    to_slogic(132),
    to_slogic(144),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(149),
    to_slogic(101),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(101),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(92),
    to_slogic(100),
    to_slogic(124),
    to_slogic(143),
    to_slogic(152),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(144),
    to_slogic(121),
    to_slogic(102),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(82),
    to_slogic(102),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(92),
    to_slogic(102),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(115),
    to_slogic(99),
    to_slogic(92),
    to_slogic(178),
    to_slogic(222),
    to_slogic(213),
    to_slogic(205),
    to_slogic(151),
    to_slogic(100),
    to_slogic(100),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(119),
    to_slogic(119),
    to_slogic(109),
    to_slogic(124),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(126),
    to_slogic(119),
    to_slogic(128),
    to_slogic(103),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(71),
    to_slogic(64),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(75),
    to_slogic(82),
    to_slogic(69),
    to_slogic(83),
    to_slogic(63),
    to_slogic(50),
    to_slogic(83),
    to_slogic(36),
    to_slogic(58),
    to_slogic(97),
    to_slogic(130),
    to_slogic(84),
    to_slogic(75),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(36),
    to_slogic(40),
    to_slogic(49),
    to_slogic(120),
    to_slogic(126),
    to_slogic(96),
    to_slogic(117),
    to_slogic(170),
    to_slogic(134),
    to_slogic(152),
    to_slogic(170),
    to_slogic(182),
    to_slogic(182),
    to_slogic(189),
    to_slogic(191),
    to_slogic(189),
    to_slogic(176),
    to_slogic(176),
    to_slogic(158),
    to_slogic(165),
    to_slogic(167),
    to_slogic(170),
    to_slogic(177),
    to_slogic(182),
    to_slogic(172),
    to_slogic(165),
    to_slogic(169),
    to_slogic(172),
    to_slogic(187),
    to_slogic(187),
    to_slogic(195),
    to_slogic(193),
    to_slogic(200),
    to_slogic(195),
    to_slogic(200),
    to_slogic(195),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(193),
    to_slogic(172),
    to_slogic(139),
    to_slogic(99),
    to_slogic(82),
    to_slogic(44),
    to_slogic(46),
    to_slogic(49),
    to_slogic(81),
    to_slogic(75),
    to_slogic(126),
    to_slogic(134),
    to_slogic(155),
    to_slogic(149),
    to_slogic(82),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(50),
    to_slogic(87),
    to_slogic(125),
    to_slogic(139),
    to_slogic(139),
    to_slogic(125),
    to_slogic(141),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(156),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(162),
    to_slogic(150),
    to_slogic(155),
    to_slogic(151),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(96),
    to_slogic(100),
    to_slogic(92),
    to_slogic(89),
    to_slogic(100),
    to_slogic(130),
    to_slogic(135),
    to_slogic(152),
    to_slogic(157),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(165),
    to_slogic(157),
    to_slogic(144),
    to_slogic(130),
    to_slogic(100),
    to_slogic(81),
    to_slogic(63),
    to_slogic(76),
    to_slogic(81),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(99),
    to_slogic(152),
    to_slogic(213),
    to_slogic(213),
    to_slogic(197),
    to_slogic(121),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(119),
    to_slogic(110),
    to_slogic(117),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(110),
    to_slogic(119),
    to_slogic(110),
    to_slogic(119),
    to_slogic(110),
    to_slogic(101),
    to_slogic(56),
    to_slogic(44),
    to_slogic(69),
    to_slogic(87),
    to_slogic(40),
    to_slogic(44),
    to_slogic(46),
    to_slogic(49),
    to_slogic(46),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(69),
    to_slogic(69),
    to_slogic(75),
    to_slogic(56),
    to_slogic(84),
    to_slogic(49),
    to_slogic(56),
    to_slogic(65),
    to_slogic(130),
    to_slogic(75),
    to_slogic(71),
    to_slogic(71),
    to_slogic(40),
    to_slogic(33),
    to_slogic(33),
    to_slogic(42),
    to_slogic(114),
    to_slogic(152),
    to_slogic(110),
    to_slogic(126),
    to_slogic(171),
    to_slogic(162),
    to_slogic(155),
    to_slogic(130),
    to_slogic(179),
    to_slogic(177),
    to_slogic(176),
    to_slogic(191),
    to_slogic(185),
    to_slogic(185),
    to_slogic(172),
    to_slogic(158),
    to_slogic(158),
    to_slogic(158),
    to_slogic(165),
    to_slogic(185),
    to_slogic(182),
    to_slogic(165),
    to_slogic(155),
    to_slogic(165),
    to_slogic(172),
    to_slogic(187),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(195),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(211),
    to_slogic(204),
    to_slogic(204),
    to_slogic(200),
    to_slogic(177),
    to_slogic(149),
    to_slogic(99),
    to_slogic(82),
    to_slogic(56),
    to_slogic(44),
    to_slogic(46),
    to_slogic(69),
    to_slogic(69),
    to_slogic(109),
    to_slogic(155),
    to_slogic(162),
    to_slogic(144),
    to_slogic(69),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(69),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(109),
    to_slogic(139),
    to_slogic(139),
    to_slogic(125),
    to_slogic(139),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(158),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(109),
    to_slogic(121),
    to_slogic(143),
    to_slogic(152),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(156),
    to_slogic(144),
    to_slogic(130),
    to_slogic(102),
    to_slogic(82),
    to_slogic(70),
    to_slogic(81),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(128),
    to_slogic(116),
    to_slogic(115),
    to_slogic(116),
    to_slogic(109),
    to_slogic(115),
    to_slogic(102),
    to_slogic(99),
    to_slogic(124),
    to_slogic(213),
    to_slogic(213),
    to_slogic(177),
    to_slogic(115),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(110),
    to_slogic(133),
    to_slogic(128),
    to_slogic(119),
    to_slogic(126),
    to_slogic(102),
    to_slogic(83),
    to_slogic(96),
    to_slogic(82),
    to_slogic(69),
    to_slogic(75),
    to_slogic(64),
    to_slogic(46),
    to_slogic(89),
    to_slogic(69),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(65),
    to_slogic(63),
    to_slogic(69),
    to_slogic(84),
    to_slogic(50),
    to_slogic(65),
    to_slogic(58),
    to_slogic(127),
    to_slogic(63),
    to_slogic(40),
    to_slogic(40),
    to_slogic(33),
    to_slogic(33),
    to_slogic(36),
    to_slogic(109),
    to_slogic(150),
    to_slogic(110),
    to_slogic(133),
    to_slogic(176),
    to_slogic(171),
    to_slogic(162),
    to_slogic(149),
    to_slogic(136),
    to_slogic(162),
    to_slogic(166),
    to_slogic(172),
    to_slogic(189),
    to_slogic(182),
    to_slogic(182),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(176),
    to_slogic(176),
    to_slogic(152),
    to_slogic(157),
    to_slogic(162),
    to_slogic(172),
    to_slogic(172),
    to_slogic(179),
    to_slogic(187),
    to_slogic(193),
    to_slogic(200),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(211),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(187),
    to_slogic(157),
    to_slogic(115),
    to_slogic(97),
    to_slogic(62),
    to_slogic(36),
    to_slogic(44),
    to_slogic(49),
    to_slogic(75),
    to_slogic(81),
    to_slogic(148),
    to_slogic(162),
    to_slogic(157),
    to_slogic(69),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(83),
    to_slogic(125),
    to_slogic(141),
    to_slogic(139),
    to_slogic(125),
    to_slogic(144),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(166),
    to_slogic(158),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(151),
    to_slogic(149),
    to_slogic(102),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(92),
    to_slogic(89),
    to_slogic(100),
    to_slogic(130),
    to_slogic(139),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(165),
    to_slogic(157),
    to_slogic(143),
    to_slogic(130),
    to_slogic(102),
    to_slogic(82),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(89),
    to_slogic(89),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(102),
    to_slogic(99),
    to_slogic(99),
    to_slogic(102),
    to_slogic(133),
    to_slogic(152),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(183),
    to_slogic(223),
    to_slogic(165),
    to_slogic(116),
    to_slogic(115),
    to_slogic(117),
    to_slogic(117),
    to_slogic(102),
    to_slogic(102),
    to_slogic(128),
    to_slogic(134),
    to_slogic(128),
    to_slogic(127),
    to_slogic(96),
    to_slogic(101),
    to_slogic(81),
    to_slogic(75),
    to_slogic(69),
    to_slogic(56),
    to_slogic(69),
    to_slogic(50),
    to_slogic(46),
    to_slogic(102),
    to_slogic(56),
    to_slogic(42),
    to_slogic(46),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(91),
    to_slogic(88),
    to_slogic(76),
    to_slogic(50),
    to_slogic(102),
    to_slogic(83),
    to_slogic(40),
    to_slogic(36),
    to_slogic(36),
    to_slogic(36),
    to_slogic(91),
    to_slogic(149),
    to_slogic(128),
    to_slogic(127),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(138),
    to_slogic(170),
    to_slogic(170),
    to_slogic(170),
    to_slogic(191),
    to_slogic(185),
    to_slogic(170),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(172),
    to_slogic(187),
    to_slogic(187),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(211),
    to_slogic(200),
    to_slogic(211),
    to_slogic(204),
    to_slogic(204),
    to_slogic(193),
    to_slogic(172),
    to_slogic(126),
    to_slogic(99),
    to_slogic(62),
    to_slogic(46),
    to_slogic(44),
    to_slogic(44),
    to_slogic(64),
    to_slogic(64),
    to_slogic(133),
    to_slogic(155),
    to_slogic(158),
    to_slogic(87),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(96),
    to_slogic(132),
    to_slogic(143),
    to_slogic(137),
    to_slogic(132),
    to_slogic(155),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(149),
    to_slogic(155),
    to_slogic(151),
    to_slogic(149),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(166),
    to_slogic(156),
    to_slogic(158),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(151),
    to_slogic(102),
    to_slogic(109),
    to_slogic(101),
    to_slogic(109),
    to_slogic(102),
    to_slogic(96),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(92),
    to_slogic(92),
    to_slogic(109),
    to_slogic(121),
    to_slogic(143),
    to_slogic(152),
    to_slogic(157),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(144),
    to_slogic(126),
    to_slogic(109),
    to_slogic(82),
    to_slogic(70),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(99),
    to_slogic(102),
    to_slogic(99),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(115),
    to_slogic(130),
    to_slogic(116),
    to_slogic(115),
    to_slogic(117),
    to_slogic(116),
    to_slogic(115),
    to_slogic(117),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(135),
    to_slogic(223),
    to_slogic(178),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(109),
    to_slogic(117),
    to_slogic(126),
    to_slogic(119),
    to_slogic(128),
    to_slogic(128),
    to_slogic(142),
    to_slogic(119),
    to_slogic(103),
    to_slogic(103),
    to_slogic(75),
    to_slogic(64),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(50),
    to_slogic(95),
    to_slogic(46),
    to_slogic(46),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(50),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(49),
    to_slogic(63),
    to_slogic(50),
    to_slogic(56),
    to_slogic(84),
    to_slogic(102),
    to_slogic(97),
    to_slogic(58),
    to_slogic(75),
    to_slogic(115),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(87),
    to_slogic(150),
    to_slogic(128),
    to_slogic(127),
    to_slogic(172),
    to_slogic(172),
    to_slogic(182),
    to_slogic(176),
    to_slogic(172),
    to_slogic(171),
    to_slogic(138),
    to_slogic(165),
    to_slogic(167),
    to_slogic(185),
    to_slogic(196),
    to_slogic(189),
    to_slogic(172),
    to_slogic(170),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(149),
    to_slogic(157),
    to_slogic(165),
    to_slogic(169),
    to_slogic(172),
    to_slogic(187),
    to_slogic(193),
    to_slogic(187),
    to_slogic(193),
    to_slogic(200),
    to_slogic(195),
    to_slogic(200),
    to_slogic(204),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(204),
    to_slogic(211),
    to_slogic(204),
    to_slogic(193),
    to_slogic(177),
    to_slogic(139),
    to_slogic(97),
    to_slogic(76),
    to_slogic(44),
    to_slogic(33),
    to_slogic(36),
    to_slogic(49),
    to_slogic(75),
    to_slogic(110),
    to_slogic(162),
    to_slogic(158),
    to_slogic(96),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(63),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(64),
    to_slogic(109),
    to_slogic(139),
    to_slogic(139),
    to_slogic(125),
    to_slogic(143),
    to_slogic(156),
    to_slogic(166),
    to_slogic(158),
    to_slogic(158),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(166),
    to_slogic(156),
    to_slogic(165),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(143),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(102),
    to_slogic(94),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(100),
    to_slogic(121),
    to_slogic(135),
    to_slogic(151),
    to_slogic(157),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(157),
    to_slogic(143),
    to_slogic(130),
    to_slogic(102),
    to_slogic(83),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(87),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(102),
    to_slogic(102),
    to_slogic(99),
    to_slogic(115),
    to_slogic(117),
    to_slogic(115),
    to_slogic(109),
    to_slogic(116),
    to_slogic(118),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(115),
    to_slogic(109),
    to_slogic(109),
    to_slogic(191),
    to_slogic(198),
    to_slogic(121),
    to_slogic(116),
    to_slogic(115),
    to_slogic(109),
    to_slogic(126),
    to_slogic(126),
    to_slogic(128),
    to_slogic(119),
    to_slogic(134),
    to_slogic(126),
    to_slogic(102),
    to_slogic(102),
    to_slogic(64),
    to_slogic(50),
    to_slogic(56),
    to_slogic(63),
    to_slogic(46),
    to_slogic(40),
    to_slogic(42),
    to_slogic(89),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(50),
    to_slogic(49),
    to_slogic(64),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(42),
    to_slogic(65),
    to_slogic(84),
    to_slogic(82),
    to_slogic(84),
    to_slogic(78),
    to_slogic(84),
    to_slogic(138),
    to_slogic(56),
    to_slogic(36),
    to_slogic(68),
    to_slogic(139),
    to_slogic(130),
    to_slogic(120),
    to_slogic(162),
    to_slogic(176),
    to_slogic(172),
    to_slogic(182),
    to_slogic(182),
    to_slogic(176),
    to_slogic(170),
    to_slogic(148),
    to_slogic(162),
    to_slogic(165),
    to_slogic(185),
    to_slogic(196),
    to_slogic(185),
    to_slogic(165),
    to_slogic(167),
    to_slogic(162),
    to_slogic(162),
    to_slogic(151),
    to_slogic(151),
    to_slogic(162),
    to_slogic(162),
    to_slogic(165),
    to_slogic(172),
    to_slogic(177),
    to_slogic(179),
    to_slogic(193),
    to_slogic(193),
    to_slogic(195),
    to_slogic(195),
    to_slogic(198),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(200),
    to_slogic(187),
    to_slogic(144),
    to_slogic(99),
    to_slogic(89),
    to_slogic(56),
    to_slogic(36),
    to_slogic(40),
    to_slogic(44),
    to_slogic(75),
    to_slogic(96),
    to_slogic(171),
    to_slogic(158),
    to_slogic(96),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(69),
    to_slogic(64),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(87),
    to_slogic(132),
    to_slogic(143),
    to_slogic(139),
    to_slogic(130),
    to_slogic(151),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(157),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(157),
    to_slogic(151),
    to_slogic(152),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(92),
    to_slogic(100),
    to_slogic(97),
    to_slogic(92),
    to_slogic(99),
    to_slogic(89),
    to_slogic(100),
    to_slogic(124),
    to_slogic(135),
    to_slogic(152),
    to_slogic(157),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(176),
    to_slogic(173),
    to_slogic(172),
    to_slogic(165),
    to_slogic(152),
    to_slogic(144),
    to_slogic(130),
    to_slogic(102),
    to_slogic(82),
    to_slogic(75),
    to_slogic(82),
    to_slogic(87),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(99),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(128),
    to_slogic(116),
    to_slogic(115),
    to_slogic(117),
    to_slogic(121),
    to_slogic(118),
    to_slogic(117),
    to_slogic(124),
    to_slogic(117),
    to_slogic(115),
    to_slogic(117),
    to_slogic(143),
    to_slogic(197),
    to_slogic(135),
    to_slogic(116),
    to_slogic(102),
    to_slogic(126),
    to_slogic(133),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(128),
    to_slogic(109),
    to_slogic(82),
    to_slogic(63),
    to_slogic(50),
    to_slogic(64),
    to_slogic(91),
    to_slogic(63),
    to_slogic(40),
    to_slogic(40),
    to_slogic(46),
    to_slogic(63),
    to_slogic(88),
    to_slogic(56),
    to_slogic(49),
    to_slogic(65),
    to_slogic(63),
    to_slogic(44),
    to_slogic(50),
    to_slogic(50),
    to_slogic(49),
    to_slogic(65),
    to_slogic(56),
    to_slogic(46),
    to_slogic(56),
    to_slogic(76),
    to_slogic(75),
    to_slogic(65),
    to_slogic(42),
    to_slogic(42),
    to_slogic(120),
    to_slogic(58),
    to_slogic(56),
    to_slogic(130),
    to_slogic(133),
    to_slogic(127),
    to_slogic(152),
    to_slogic(173),
    to_slogic(166),
    to_slogic(177),
    to_slogic(189),
    to_slogic(185),
    to_slogic(185),
    to_slogic(165),
    to_slogic(143),
    to_slogic(153),
    to_slogic(176),
    to_slogic(191),
    to_slogic(191),
    to_slogic(176),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(169),
    to_slogic(172),
    to_slogic(187),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(195),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(214),
    to_slogic(200),
    to_slogic(193),
    to_slogic(151),
    to_slogic(118),
    to_slogic(89),
    to_slogic(56),
    to_slogic(46),
    to_slogic(40),
    to_slogic(46),
    to_slogic(63),
    to_slogic(75),
    to_slogic(162),
    to_slogic(162),
    to_slogic(109),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(109),
    to_slogic(141),
    to_slogic(139),
    to_slogic(132),
    to_slogic(139),
    to_slogic(156),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(156),
    to_slogic(166),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(149),
    to_slogic(156),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(143),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(101),
    to_slogic(100),
    to_slogic(102),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(100),
    to_slogic(130),
    to_slogic(135),
    to_slogic(152),
    to_slogic(157),
    to_slogic(173),
    to_slogic(165),
    to_slogic(176),
    to_slogic(172),
    to_slogic(178),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(157),
    to_slogic(151),
    to_slogic(130),
    to_slogic(102),
    to_slogic(75),
    to_slogic(77),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(99),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(117),
    to_slogic(121),
    to_slogic(116),
    to_slogic(121),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(116),
    to_slogic(124),
    to_slogic(126),
    to_slogic(151),
    to_slogic(121),
    to_slogic(116),
    to_slogic(121),
    to_slogic(139),
    to_slogic(134),
    to_slogic(133),
    to_slogic(128),
    to_slogic(128),
    to_slogic(117),
    to_slogic(82),
    to_slogic(49),
    to_slogic(63),
    to_slogic(50),
    to_slogic(42),
    to_slogic(89),
    to_slogic(50),
    to_slogic(46),
    to_slogic(56),
    to_slogic(46),
    to_slogic(46),
    to_slogic(75),
    to_slogic(56),
    to_slogic(56),
    to_slogic(81),
    to_slogic(56),
    to_slogic(46),
    to_slogic(49),
    to_slogic(46),
    to_slogic(50),
    to_slogic(75),
    to_slogic(69),
    to_slogic(50),
    to_slogic(46),
    to_slogic(56),
    to_slogic(65),
    to_slogic(71),
    to_slogic(36),
    to_slogic(36),
    to_slogic(81),
    to_slogic(97),
    to_slogic(120),
    to_slogic(137),
    to_slogic(117),
    to_slogic(141),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(176),
    to_slogic(182),
    to_slogic(185),
    to_slogic(191),
    to_slogic(170),
    to_slogic(143),
    to_slogic(148),
    to_slogic(185),
    to_slogic(189),
    to_slogic(172),
    to_slogic(158),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(157),
    to_slogic(161),
    to_slogic(162),
    to_slogic(169),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(177),
    to_slogic(176),
    to_slogic(187),
    to_slogic(195),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(204),
    to_slogic(195),
    to_slogic(162),
    to_slogic(124),
    to_slogic(99),
    to_slogic(76),
    to_slogic(49),
    to_slogic(46),
    to_slogic(40),
    to_slogic(50),
    to_slogic(81),
    to_slogic(144),
    to_slogic(171),
    to_slogic(101),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(75),
    to_slogic(120),
    to_slogic(143),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(156),
    to_slogic(166),
    to_slogic(156),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(166),
    to_slogic(166),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(152),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(89),
    to_slogic(102),
    to_slogic(116),
    to_slogic(143),
    to_slogic(144),
    to_slogic(157),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(176),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(144),
    to_slogic(130),
    to_slogic(100),
    to_slogic(81),
    to_slogic(77),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(115),
    to_slogic(102),
    to_slogic(109),
    to_slogic(121),
    to_slogic(116),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(100),
    to_slogic(121),
    to_slogic(136),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(115),
    to_slogic(130),
    to_slogic(124),
    to_slogic(133),
    to_slogic(133),
    to_slogic(122),
    to_slogic(121),
    to_slogic(96),
    to_slogic(69),
    to_slogic(50),
    to_slogic(71),
    to_slogic(42),
    to_slogic(42),
    to_slogic(97),
    to_slogic(56),
    to_slogic(65),
    to_slogic(49),
    to_slogic(50),
    to_slogic(36),
    to_slogic(49),
    to_slogic(69),
    to_slogic(89),
    to_slogic(75),
    to_slogic(44),
    to_slogic(44),
    to_slogic(50),
    to_slogic(46),
    to_slogic(63),
    to_slogic(69),
    to_slogic(50),
    to_slogic(69),
    to_slogic(50),
    to_slogic(50),
    to_slogic(71),
    to_slogic(95),
    to_slogic(33),
    to_slogic(33),
    to_slogic(40),
    to_slogic(110),
    to_slogic(139),
    to_slogic(119),
    to_slogic(141),
    to_slogic(172),
    to_slogic(162),
    to_slogic(162),
    to_slogic(157),
    to_slogic(167),
    to_slogic(185),
    to_slogic(189),
    to_slogic(185),
    to_slogic(177),
    to_slogic(162),
    to_slogic(165),
    to_slogic(177),
    to_slogic(176),
    to_slogic(162),
    to_slogic(162),
    to_slogic(151),
    to_slogic(161),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(169),
    to_slogic(172),
    to_slogic(169),
    to_slogic(187),
    to_slogic(172),
    to_slogic(187),
    to_slogic(187),
    to_slogic(195),
    to_slogic(195),
    to_slogic(193),
    to_slogic(195),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(198),
    to_slogic(172),
    to_slogic(134),
    to_slogic(99),
    to_slogic(81),
    to_slogic(46),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(81),
    to_slogic(132),
    to_slogic(172),
    to_slogic(120),
    to_slogic(64),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(63),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(95),
    to_slogic(132),
    to_slogic(139),
    to_slogic(130),
    to_slogic(139),
    to_slogic(150),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(156),
    to_slogic(166),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(166),
    to_slogic(156),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(149),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(143),
    to_slogic(151),
    to_slogic(102),
    to_slogic(109),
    to_slogic(94),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(100),
    to_slogic(94),
    to_slogic(89),
    to_slogic(89),
    to_slogic(100),
    to_slogic(124),
    to_slogic(139),
    to_slogic(152),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(156),
    to_slogic(143),
    to_slogic(130),
    to_slogic(100),
    to_slogic(82),
    to_slogic(70),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(96),
    to_slogic(99),
    to_slogic(102),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(99),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(115),
    to_slogic(124),
    to_slogic(116),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(116),
    to_slogic(133),
    to_slogic(117),
    to_slogic(101),
    to_slogic(137),
    to_slogic(150),
    to_slogic(118),
    to_slogic(119),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(119),
    to_slogic(119),
    to_slogic(92),
    to_slogic(50),
    to_slogic(76),
    to_slogic(83),
    to_slogic(36),
    to_slogic(42),
    to_slogic(102),
    to_slogic(71),
    to_slogic(50),
    to_slogic(46),
    to_slogic(49),
    to_slogic(63),
    to_slogic(69),
    to_slogic(97),
    to_slogic(75),
    to_slogic(56),
    to_slogic(44),
    to_slogic(46),
    to_slogic(50),
    to_slogic(44),
    to_slogic(75),
    to_slogic(50),
    to_slogic(50),
    to_slogic(91),
    to_slogic(50),
    to_slogic(50),
    to_slogic(89),
    to_slogic(49),
    to_slogic(42),
    to_slogic(36),
    to_slogic(81),
    to_slogic(125),
    to_slogic(96),
    to_slogic(120),
    to_slogic(176),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(167),
    to_slogic(185),
    to_slogic(191),
    to_slogic(185),
    to_slogic(185),
    to_slogic(170),
    to_slogic(177),
    to_slogic(176),
    to_slogic(167),
    to_slogic(149),
    to_slogic(151),
    to_slogic(165),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(169),
    to_slogic(169),
    to_slogic(177),
    to_slogic(169),
    to_slogic(176),
    to_slogic(172),
    to_slogic(172),
    to_slogic(187),
    to_slogic(179),
    to_slogic(193),
    to_slogic(195),
    to_slogic(193),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(187),
    to_slogic(139),
    to_slogic(99),
    to_slogic(81),
    to_slogic(56),
    to_slogic(36),
    to_slogic(44),
    to_slogic(46),
    to_slogic(75),
    to_slogic(110),
    to_slogic(176),
    to_slogic(126),
    to_slogic(69),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(63),
    to_slogic(120),
    to_slogic(141),
    to_slogic(139),
    to_slogic(125),
    to_slogic(139),
    to_slogic(156),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(158),
    to_slogic(162),
    to_slogic(166),
    to_slogic(158),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(158),
    to_slogic(166),
    to_slogic(158),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(132),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(143),
    to_slogic(155),
    to_slogic(155),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(92),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(89),
    to_slogic(102),
    to_slogic(124),
    to_slogic(144),
    to_slogic(152),
    to_slogic(157),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(176),
    to_slogic(173),
    to_slogic(165),
    to_slogic(165),
    to_slogic(143),
    to_slogic(130),
    to_slogic(100),
    to_slogic(82),
    to_slogic(77),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(115),
    to_slogic(115),
    to_slogic(109),
    to_slogic(116),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(117),
    to_slogic(121),
    to_slogic(128),
    to_slogic(143),
    to_slogic(144),
    to_slogic(109),
    to_slogic(121),
    to_slogic(161),
    to_slogic(134),
    to_slogic(121),
    to_slogic(122),
    to_slogic(134),
    to_slogic(119),
    to_slogic(119),
    to_slogic(110),
    to_slogic(64),
    to_slogic(58),
    to_slogic(89),
    to_slogic(65),
    to_slogic(36),
    to_slogic(50),
    to_slogic(107),
    to_slogic(75),
    to_slogic(36),
    to_slogic(49),
    to_slogic(46),
    to_slogic(75),
    to_slogic(89),
    to_slogic(75),
    to_slogic(63),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(50),
    to_slogic(49),
    to_slogic(83),
    to_slogic(40),
    to_slogic(42),
    to_slogic(97),
    to_slogic(50),
    to_slogic(63),
    to_slogic(71),
    to_slogic(50),
    to_slogic(50),
    to_slogic(64),
    to_slogic(139),
    to_slogic(117),
    to_slogic(110),
    to_slogic(182),
    to_slogic(173),
    to_slogic(166),
    to_slogic(176),
    to_slogic(167),
    to_slogic(156),
    to_slogic(165),
    to_slogic(185),
    to_slogic(191),
    to_slogic(191),
    to_slogic(185),
    to_slogic(177),
    to_slogic(176),
    to_slogic(137),
    to_slogic(117),
    to_slogic(128),
    to_slogic(146),
    to_slogic(149),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(169),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(177),
    to_slogic(172),
    to_slogic(177),
    to_slogic(187),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(195),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(198),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(204),
    to_slogic(198),
    to_slogic(177),
    to_slogic(146),
    to_slogic(99),
    to_slogic(56),
    to_slogic(56),
    to_slogic(36),
    to_slogic(44),
    to_slogic(46),
    to_slogic(69),
    to_slogic(95),
    to_slogic(176),
    to_slogic(141),
    to_slogic(69),
    to_slogic(69),
    to_slogic(56),
    to_slogic(68),
    to_slogic(63),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(87),
    to_slogic(120),
    to_slogic(139),
    to_slogic(130),
    to_slogic(134),
    to_slogic(143),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(166),
    to_slogic(166),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(121),
    to_slogic(139),
    to_slogic(152),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(172),
    to_slogic(157),
    to_slogic(143),
    to_slogic(130),
    to_slogic(100),
    to_slogic(82),
    to_slogic(76),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(99),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(121),
    to_slogic(115),
    to_slogic(116),
    to_slogic(121),
    to_slogic(116),
    to_slogic(121),
    to_slogic(118),
    to_slogic(172),
    to_slogic(178),
    to_slogic(136),
    to_slogic(76),
    to_slogic(40),
    to_slogic(44),
    to_slogic(62),
    to_slogic(121),
    to_slogic(141),
    to_slogic(133),
    to_slogic(124),
    to_slogic(109),
    to_slogic(109),
    to_slogic(77),
    to_slogic(56),
    to_slogic(78),
    to_slogic(97),
    to_slogic(42),
    to_slogic(42),
    to_slogic(65),
    to_slogic(120),
    to_slogic(50),
    to_slogic(33),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(42),
    to_slogic(49),
    to_slogic(46),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(42),
    to_slogic(65),
    to_slogic(97),
    to_slogic(46),
    to_slogic(76),
    to_slogic(56),
    to_slogic(42),
    to_slogic(49),
    to_slogic(120),
    to_slogic(133),
    to_slogic(101),
    to_slogic(162),
    to_slogic(177),
    to_slogic(166),
    to_slogic(177),
    to_slogic(182),
    to_slogic(166),
    to_slogic(151),
    to_slogic(162),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(171),
    to_slogic(118),
    to_slogic(81),
    to_slogic(92),
    to_slogic(102),
    to_slogic(109),
    to_slogic(119),
    to_slogic(119),
    to_slogic(134),
    to_slogic(149),
    to_slogic(155),
    to_slogic(169),
    to_slogic(169),
    to_slogic(177),
    to_slogic(176),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(177),
    to_slogic(187),
    to_slogic(193),
    to_slogic(195),
    to_slogic(193),
    to_slogic(187),
    to_slogic(195),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(207),
    to_slogic(204),
    to_slogic(200),
    to_slogic(187),
    to_slogic(162),
    to_slogic(130),
    to_slogic(76),
    to_slogic(56),
    to_slogic(44),
    to_slogic(33),
    to_slogic(44),
    to_slogic(36),
    to_slogic(75),
    to_slogic(81),
    to_slogic(176),
    to_slogic(149),
    to_slogic(83),
    to_slogic(56),
    to_slogic(69),
    to_slogic(63),
    to_slogic(64),
    to_slogic(56),
    to_slogic(63),
    to_slogic(68),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(101),
    to_slogic(132),
    to_slogic(139),
    to_slogic(134),
    to_slogic(132),
    to_slogic(149),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(158),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(166),
    to_slogic(162),
    to_slogic(166),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(143),
    to_slogic(133),
    to_slogic(139),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(96),
    to_slogic(102),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(121),
    to_slogic(139),
    to_slogic(152),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(178),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(144),
    to_slogic(130),
    to_slogic(100),
    to_slogic(75),
    to_slogic(77),
    to_slogic(83),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(115),
    to_slogic(117),
    to_slogic(121),
    to_slogic(117),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(183),
    to_slogic(144),
    to_slogic(70),
    to_slogic(44),
    to_slogic(36),
    to_slogic(44),
    to_slogic(81),
    to_slogic(148),
    to_slogic(193),
    to_slogic(162),
    to_slogic(102),
    to_slogic(89),
    to_slogic(82),
    to_slogic(50),
    to_slogic(65),
    to_slogic(89),
    to_slogic(89),
    to_slogic(42),
    to_slogic(44),
    to_slogic(89),
    to_slogic(130),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(64),
    to_slogic(84),
    to_slogic(64),
    to_slogic(65),
    to_slogic(75),
    to_slogic(56),
    to_slogic(65),
    to_slogic(42),
    to_slogic(40),
    to_slogic(96),
    to_slogic(137),
    to_slogic(96),
    to_slogic(144),
    to_slogic(177),
    to_slogic(166),
    to_slogic(183),
    to_slogic(189),
    to_slogic(182),
    to_slogic(162),
    to_slogic(157),
    to_slogic(176),
    to_slogic(185),
    to_slogic(196),
    to_slogic(189),
    to_slogic(171),
    to_slogic(128),
    to_slogic(119),
    to_slogic(128),
    to_slogic(127),
    to_slogic(118),
    to_slogic(101),
    to_slogic(92),
    to_slogic(82),
    to_slogic(82),
    to_slogic(99),
    to_slogic(119),
    to_slogic(146),
    to_slogic(165),
    to_slogic(172),
    to_slogic(177),
    to_slogic(172),
    to_slogic(169),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(187),
    to_slogic(187),
    to_slogic(193),
    to_slogic(187),
    to_slogic(187),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(198),
    to_slogic(200),
    to_slogic(200),
    to_slogic(193),
    to_slogic(177),
    to_slogic(152),
    to_slogic(128),
    to_slogic(102),
    to_slogic(63),
    to_slogic(56),
    to_slogic(44),
    to_slogic(36),
    to_slogic(40),
    to_slogic(44),
    to_slogic(68),
    to_slogic(69),
    to_slogic(165),
    to_slogic(157),
    to_slogic(96),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(69),
    to_slogic(110),
    to_slogic(139),
    to_slogic(141),
    to_slogic(125),
    to_slogic(139),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(158),
    to_slogic(149),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(132),
    to_slogic(144),
    to_slogic(141),
    to_slogic(133),
    to_slogic(139),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(124),
    to_slogic(144),
    to_slogic(144),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(157),
    to_slogic(143),
    to_slogic(135),
    to_slogic(100),
    to_slogic(82),
    to_slogic(77),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(99),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(119),
    to_slogic(134),
    to_slogic(133),
    to_slogic(151),
    to_slogic(157),
    to_slogic(94),
    to_slogic(62),
    to_slogic(40),
    to_slogic(42),
    to_slogic(96),
    to_slogic(151),
    to_slogic(128),
    to_slogic(109),
    to_slogic(82),
    to_slogic(69),
    to_slogic(75),
    to_slogic(63),
    to_slogic(78),
    to_slogic(97),
    to_slogic(50),
    to_slogic(42),
    to_slogic(76),
    to_slogic(84),
    to_slogic(113),
    to_slogic(56),
    to_slogic(36),
    to_slogic(42),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(75),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(36),
    to_slogic(75),
    to_slogic(76),
    to_slogic(89),
    to_slogic(56),
    to_slogic(65),
    to_slogic(56),
    to_slogic(36),
    to_slogic(68),
    to_slogic(144),
    to_slogic(117),
    to_slogic(141),
    to_slogic(176),
    to_slogic(162),
    to_slogic(183),
    to_slogic(182),
    to_slogic(196),
    to_slogic(171),
    to_slogic(149),
    to_slogic(162),
    to_slogic(185),
    to_slogic(191),
    to_slogic(196),
    to_slogic(156),
    to_slogic(126),
    to_slogic(139),
    to_slogic(146),
    to_slogic(151),
    to_slogic(149),
    to_slogic(151),
    to_slogic(149),
    to_slogic(126),
    to_slogic(92),
    to_slogic(76),
    to_slogic(63),
    to_slogic(62),
    to_slogic(81),
    to_slogic(109),
    to_slogic(149),
    to_slogic(162),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(187),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(187),
    to_slogic(187),
    to_slogic(193),
    to_slogic(187),
    to_slogic(193),
    to_slogic(187),
    to_slogic(177),
    to_slogic(158),
    to_slogic(133),
    to_slogic(101),
    to_slogic(92),
    to_slogic(82),
    to_slogic(92),
    to_slogic(81),
    to_slogic(76),
    to_slogic(56),
    to_slogic(44),
    to_slogic(40),
    to_slogic(46),
    to_slogic(64),
    to_slogic(64),
    to_slogic(162),
    to_slogic(158),
    to_slogic(120),
    to_slogic(56),
    to_slogic(56),
    to_slogic(69),
    to_slogic(75),
    to_slogic(64),
    to_slogic(69),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(81),
    to_slogic(125),
    to_slogic(139),
    to_slogic(132),
    to_slogic(134),
    to_slogic(143),
    to_slogic(162),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(156),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(162),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(158),
    to_slogic(156),
    to_slogic(149),
    to_slogic(156),
    to_slogic(156),
    to_slogic(158),
    to_slogic(155),
    to_slogic(149),
    to_slogic(157),
    to_slogic(144),
    to_slogic(149),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(133),
    to_slogic(132),
    to_slogic(132),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(89),
    to_slogic(99),
    to_slogic(124),
    to_slogic(135),
    to_slogic(152),
    to_slogic(152),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(172),
    to_slogic(178),
    to_slogic(173),
    to_slogic(172),
    to_slogic(157),
    to_slogic(144),
    to_slogic(130),
    to_slogic(100),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(115),
    to_slogic(116),
    to_slogic(118),
    to_slogic(133),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(83),
    to_slogic(63),
    to_slogic(68),
    to_slogic(42),
    to_slogic(89),
    to_slogic(134),
    to_slogic(109),
    to_slogic(75),
    to_slogic(87),
    to_slogic(69),
    to_slogic(64),
    to_slogic(69),
    to_slogic(97),
    to_slogic(65),
    to_slogic(44),
    to_slogic(65),
    to_slogic(97),
    to_slogic(58),
    to_slogic(95),
    to_slogic(83),
    to_slogic(40),
    to_slogic(49),
    to_slogic(71),
    to_slogic(56),
    to_slogic(50),
    to_slogic(56),
    to_slogic(89),
    to_slogic(65),
    to_slogic(49),
    to_slogic(33),
    to_slogic(44),
    to_slogic(40),
    to_slogic(42),
    to_slogic(81),
    to_slogic(102),
    to_slogic(49),
    to_slogic(71),
    to_slogic(36),
    to_slogic(40),
    to_slogic(125),
    to_slogic(144),
    to_slogic(120),
    to_slogic(176),
    to_slogic(173),
    to_slogic(177),
    to_slogic(182),
    to_slogic(196),
    to_slogic(189),
    to_slogic(156),
    to_slogic(158),
    to_slogic(176),
    to_slogic(196),
    to_slogic(193),
    to_slogic(143),
    to_slogic(117),
    to_slogic(130),
    to_slogic(134),
    to_slogic(137),
    to_slogic(139),
    to_slogic(126),
    to_slogic(152),
    to_slogic(155),
    to_slogic(139),
    to_slogic(128),
    to_slogic(102),
    to_slogic(99),
    to_slogic(82),
    to_slogic(76),
    to_slogic(77),
    to_slogic(92),
    to_slogic(139),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(176),
    to_slogic(187),
    to_slogic(187),
    to_slogic(193),
    to_slogic(187),
    to_slogic(193),
    to_slogic(187),
    to_slogic(187),
    to_slogic(176),
    to_slogic(157),
    to_slogic(126),
    to_slogic(92),
    to_slogic(96),
    to_slogic(92),
    to_slogic(101),
    to_slogic(119),
    to_slogic(119),
    to_slogic(109),
    to_slogic(97),
    to_slogic(62),
    to_slogic(56),
    to_slogic(40),
    to_slogic(44),
    to_slogic(56),
    to_slogic(64),
    to_slogic(158),
    to_slogic(157),
    to_slogic(110),
    to_slogic(69),
    to_slogic(49),
    to_slogic(64),
    to_slogic(63),
    to_slogic(64),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(87),
    to_slogic(125),
    to_slogic(139),
    to_slogic(134),
    to_slogic(132),
    to_slogic(155),
    to_slogic(158),
    to_slogic(162),
    to_slogic(156),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(162),
    to_slogic(156),
    to_slogic(158),
    to_slogic(162),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(158),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(158),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(156),
    to_slogic(158),
    to_slogic(149),
    to_slogic(158),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(132),
    to_slogic(133),
    to_slogic(132),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(96),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(92),
    to_slogic(89),
    to_slogic(89),
    to_slogic(99),
    to_slogic(121),
    to_slogic(135),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(176),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(157),
    to_slogic(152),
    to_slogic(130),
    to_slogic(109),
    to_slogic(82),
    to_slogic(76),
    to_slogic(82),
    to_slogic(82),
    to_slogic(99),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(102),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(128),
    to_slogic(152),
    to_slogic(155),
    to_slogic(146),
    to_slogic(144),
    to_slogic(165),
    to_slogic(156),
    to_slogic(118),
    to_slogic(144),
    to_slogic(96),
    to_slogic(121),
    to_slogic(117),
    to_slogic(133),
    to_slogic(75),
    to_slogic(75),
    to_slogic(49),
    to_slogic(63),
    to_slogic(83),
    to_slogic(103),
    to_slogic(69),
    to_slogic(76),
    to_slogic(91),
    to_slogic(89),
    to_slogic(42),
    to_slogic(63),
    to_slogic(97),
    to_slogic(42),
    to_slogic(49),
    to_slogic(71),
    to_slogic(49),
    to_slogic(40),
    to_slogic(46),
    to_slogic(89),
    to_slogic(88),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(63),
    to_slogic(71),
    to_slogic(33),
    to_slogic(40),
    to_slogic(91),
    to_slogic(137),
    to_slogic(119),
    to_slogic(172),
    to_slogic(177),
    to_slogic(166),
    to_slogic(182),
    to_slogic(193),
    to_slogic(196),
    to_slogic(182),
    to_slogic(167),
    to_slogic(176),
    to_slogic(189),
    to_slogic(189),
    to_slogic(130),
    to_slogic(97),
    to_slogic(115),
    to_slogic(109),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(62),
    to_slogic(109),
    to_slogic(144),
    to_slogic(97),
    to_slogic(117),
    to_slogic(99),
    to_slogic(119),
    to_slogic(102),
    to_slogic(118),
    to_slogic(92),
    to_slogic(102),
    to_slogic(118),
    to_slogic(146),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(187),
    to_slogic(187),
    to_slogic(187),
    to_slogic(172),
    to_slogic(155),
    to_slogic(119),
    to_slogic(110),
    to_slogic(109),
    to_slogic(117),
    to_slogic(99),
    to_slogic(99),
    to_slogic(109),
    to_slogic(99),
    to_slogic(81),
    to_slogic(81),
    to_slogic(62),
    to_slogic(62),
    to_slogic(44),
    to_slogic(42),
    to_slogic(56),
    to_slogic(63),
    to_slogic(149),
    to_slogic(162),
    to_slogic(119),
    to_slogic(75),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(110),
    to_slogic(141),
    to_slogic(132),
    to_slogic(125),
    to_slogic(137),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(155),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(162),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(158),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(133),
    to_slogic(144),
    to_slogic(133),
    to_slogic(133),
    to_slogic(102),
    to_slogic(100),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(99),
    to_slogic(89),
    to_slogic(81),
    to_slogic(92),
    to_slogic(121),
    to_slogic(139),
    to_slogic(152),
    to_slogic(157),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(173),
    to_slogic(176),
    to_slogic(173),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(102),
    to_slogic(81),
    to_slogic(77),
    to_slogic(82),
    to_slogic(81),
    to_slogic(82),
    to_slogic(102),
    to_slogic(92),
    to_slogic(100),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(97),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(102),
    to_slogic(110),
    to_slogic(120),
    to_slogic(141),
    to_slogic(144),
    to_slogic(144),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(165),
    to_slogic(152),
    to_slogic(162),
    to_slogic(128),
    to_slogic(75),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(71),
    to_slogic(65),
    to_slogic(84),
    to_slogic(109),
    to_slogic(76),
    to_slogic(69),
    to_slogic(84),
    to_slogic(95),
    to_slogic(71),
    to_slogic(36),
    to_slogic(50),
    to_slogic(89),
    to_slogic(56),
    to_slogic(49),
    to_slogic(83),
    to_slogic(49),
    to_slogic(36),
    to_slogic(42),
    to_slogic(65),
    to_slogic(102),
    to_slogic(63),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(42),
    to_slogic(56),
    to_slogic(139),
    to_slogic(117),
    to_slogic(149),
    to_slogic(183),
    to_slogic(166),
    to_slogic(177),
    to_slogic(189),
    to_slogic(196),
    to_slogic(204),
    to_slogic(182),
    to_slogic(176),
    to_slogic(189),
    to_slogic(182),
    to_slogic(109),
    to_slogic(81),
    to_slogic(89),
    to_slogic(81),
    to_slogic(81),
    to_slogic(62),
    to_slogic(62),
    to_slogic(56),
    to_slogic(44),
    to_slogic(62),
    to_slogic(76),
    to_slogic(44),
    to_slogic(56),
    to_slogic(62),
    to_slogic(109),
    to_slogic(102),
    to_slogic(128),
    to_slogic(118),
    to_slogic(126),
    to_slogic(124),
    to_slogic(134),
    to_slogic(149),
    to_slogic(157),
    to_slogic(149),
    to_slogic(162),
    to_slogic(172),
    to_slogic(193),
    to_slogic(187),
    to_slogic(195),
    to_slogic(193),
    to_slogic(193),
    to_slogic(187),
    to_slogic(162),
    to_slogic(133),
    to_slogic(119),
    to_slogic(102),
    to_slogic(62),
    to_slogic(62),
    to_slogic(56),
    to_slogic(44),
    to_slogic(62),
    to_slogic(63),
    to_slogic(62),
    to_slogic(62),
    to_slogic(70),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(69),
    to_slogic(143),
    to_slogic(162),
    to_slogic(109),
    to_slogic(83),
    to_slogic(56),
    to_slogic(56),
    to_slogic(69),
    to_slogic(63),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(83),
    to_slogic(125),
    to_slogic(139),
    to_slogic(132),
    to_slogic(134),
    to_slogic(143),
    to_slogic(162),
    to_slogic(156),
    to_slogic(158),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(156),
    to_slogic(155),
    to_slogic(158),
    to_slogic(156),
    to_slogic(158),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(158),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(149),
    to_slogic(156),
    to_slogic(158),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(133),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(100),
    to_slogic(81),
    to_slogic(81),
    to_slogic(99),
    to_slogic(121),
    to_slogic(135),
    to_slogic(144),
    to_slogic(157),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(173),
    to_slogic(172),
    to_slogic(157),
    to_slogic(151),
    to_slogic(130),
    to_slogic(109),
    to_slogic(82),
    to_slogic(76),
    to_slogic(76),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(92),
    to_slogic(97),
    to_slogic(99),
    to_slogic(103),
    to_slogic(144),
    to_slogic(172),
    to_slogic(157),
    to_slogic(137),
    to_slogic(151),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(139),
    to_slogic(96),
    to_slogic(119),
    to_slogic(96),
    to_slogic(44),
    to_slogic(40),
    to_slogic(42),
    to_slogic(71),
    to_slogic(91),
    to_slogic(78),
    to_slogic(107),
    to_slogic(115),
    to_slogic(69),
    to_slogic(78),
    to_slogic(91),
    to_slogic(102),
    to_slogic(71),
    to_slogic(42),
    to_slogic(56),
    to_slogic(65),
    to_slogic(65),
    to_slogic(50),
    to_slogic(89),
    to_slogic(49),
    to_slogic(40),
    to_slogic(36),
    to_slogic(42),
    to_slogic(83),
    to_slogic(107),
    to_slogic(71),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(33),
    to_slogic(36),
    to_slogic(40),
    to_slogic(114),
    to_slogic(137),
    to_slogic(125),
    to_slogic(182),
    to_slogic(173),
    to_slogic(177),
    to_slogic(182),
    to_slogic(200),
    to_slogic(200),
    to_slogic(191),
    to_slogic(182),
    to_slogic(189),
    to_slogic(171),
    to_slogic(94),
    to_slogic(76),
    to_slogic(62),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(102),
    to_slogic(139),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(139),
    to_slogic(142),
    to_slogic(146),
    to_slogic(152),
    to_slogic(162),
    to_slogic(169),
    to_slogic(187),
    to_slogic(195),
    to_slogic(200),
    to_slogic(198),
    to_slogic(193),
    to_slogic(173),
    to_slogic(128),
    to_slogic(89),
    to_slogic(62),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(62),
    to_slogic(44),
    to_slogic(44),
    to_slogic(36),
    to_slogic(56),
    to_slogic(64),
    to_slogic(133),
    to_slogic(172),
    to_slogic(120),
    to_slogic(87),
    to_slogic(64),
    to_slogic(56),
    to_slogic(75),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(42),
    to_slogic(87),
    to_slogic(139),
    to_slogic(139),
    to_slogic(132),
    to_slogic(139),
    to_slogic(143),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(156),
    to_slogic(158),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(155),
    to_slogic(157),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(162),
    to_slogic(150),
    to_slogic(155),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(156),
    to_slogic(149),
    to_slogic(156),
    to_slogic(155),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(143),
    to_slogic(133),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(96),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(81),
    to_slogic(81),
    to_slogic(89),
    to_slogic(121),
    to_slogic(135),
    to_slogic(151),
    to_slogic(157),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(176),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(156),
    to_slogic(143),
    to_slogic(130),
    to_slogic(102),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(89),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(97),
    to_slogic(99),
    to_slogic(89),
    to_slogic(99),
    to_slogic(99),
    to_slogic(97),
    to_slogic(82),
    to_slogic(92),
    to_slogic(162),
    to_slogic(183),
    to_slogic(203),
    to_slogic(135),
    to_slogic(143),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(146),
    to_slogic(139),
    to_slogic(120),
    to_slogic(69),
    to_slogic(69),
    to_slogic(64),
    to_slogic(42),
    to_slogic(36),
    to_slogic(76),
    to_slogic(107),
    to_slogic(82),
    to_slogic(76),
    to_slogic(102),
    to_slogic(65),
    to_slogic(84),
    to_slogic(84),
    to_slogic(76),
    to_slogic(122),
    to_slogic(71),
    to_slogic(42),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(65),
    to_slogic(95),
    to_slogic(56),
    to_slogic(42),
    to_slogic(40),
    to_slogic(40),
    to_slogic(50),
    to_slogic(89),
    to_slogic(115),
    to_slogic(83),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(75),
    to_slogic(143),
    to_slogic(117),
    to_slogic(176),
    to_slogic(177),
    to_slogic(166),
    to_slogic(176),
    to_slogic(182),
    to_slogic(196),
    to_slogic(196),
    to_slogic(189),
    to_slogic(189),
    to_slogic(182),
    to_slogic(109),
    to_slogic(62),
    to_slogic(62),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(46),
    to_slogic(75),
    to_slogic(126),
    to_slogic(96),
    to_slogic(56),
    to_slogic(44),
    to_slogic(33),
    to_slogic(56),
    to_slogic(102),
    to_slogic(133),
    to_slogic(128),
    to_slogic(126),
    to_slogic(134),
    to_slogic(139),
    to_slogic(149),
    to_slogic(149),
    to_slogic(162),
    to_slogic(169),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(183),
    to_slogic(101),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(50),
    to_slogic(70),
    to_slogic(96),
    to_slogic(70),
    to_slogic(56),
    to_slogic(49),
    to_slogic(62),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(40),
    to_slogic(56),
    to_slogic(64),
    to_slogic(133),
    to_slogic(172),
    to_slogic(119),
    to_slogic(83),
    to_slogic(63),
    to_slogic(56),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(101),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(162),
    to_slogic(158),
    to_slogic(162),
    to_slogic(158),
    to_slogic(155),
    to_slogic(157),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(162),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(132),
    to_slogic(100),
    to_slogic(96),
    to_slogic(99),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(81),
    to_slogic(89),
    to_slogic(70),
    to_slogic(81),
    to_slogic(109),
    to_slogic(135),
    to_slogic(144),
    to_slogic(165),
    to_slogic(172),
    to_slogic(178),
    to_slogic(172),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(172),
    to_slogic(157),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(81),
    to_slogic(76),
    to_slogic(76),
    to_slogic(82),
    to_slogic(89),
    to_slogic(92),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(89),
    to_slogic(89),
    to_slogic(77),
    to_slogic(115),
    to_slogic(193),
    to_slogic(191),
    to_slogic(176),
    to_slogic(130),
    to_slogic(144),
    to_slogic(144),
    to_slogic(156),
    to_slogic(152),
    to_slogic(101),
    to_slogic(134),
    to_slogic(110),
    to_slogic(75),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(71),
    to_slogic(115),
    to_slogic(63),
    to_slogic(50),
    to_slogic(102),
    to_slogic(49),
    to_slogic(42),
    to_slogic(84),
    to_slogic(103),
    to_slogic(97),
    to_slogic(120),
    to_slogic(56),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(95),
    to_slogic(68),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(44),
    to_slogic(56),
    to_slogic(71),
    to_slogic(63),
    to_slogic(83),
    to_slogic(56),
    to_slogic(40),
    to_slogic(36),
    to_slogic(40),
    to_slogic(130),
    to_slogic(128),
    to_slogic(141),
    to_slogic(182),
    to_slogic(166),
    to_slogic(177),
    to_slogic(182),
    to_slogic(189),
    to_slogic(205),
    to_slogic(196),
    to_slogic(193),
    to_slogic(189),
    to_slogic(102),
    to_slogic(81),
    to_slogic(76),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(69),
    to_slogic(109),
    to_slogic(192),
    to_slogic(183),
    to_slogic(134),
    to_slogic(69),
    to_slogic(44),
    to_slogic(63),
    to_slogic(77),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(134),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(162),
    to_slogic(169),
    to_slogic(193),
    to_slogic(211),
    to_slogic(204),
    to_slogic(198),
    to_slogic(117),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(50),
    to_slogic(89),
    to_slogic(102),
    to_slogic(155),
    to_slogic(125),
    to_slogic(63),
    to_slogic(33),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(64),
    to_slogic(50),
    to_slogic(120),
    to_slogic(176),
    to_slogic(110),
    to_slogic(91),
    to_slogic(69),
    to_slogic(69),
    to_slogic(75),
    to_slogic(64),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(69),
    to_slogic(120),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(149),
    to_slogic(158),
    to_slogic(156),
    to_slogic(162),
    to_slogic(150),
    to_slogic(162),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(157),
    to_slogic(149),
    to_slogic(157),
    to_slogic(149),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(133),
    to_slogic(143),
    to_slogic(133),
    to_slogic(132),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(100),
    to_slogic(94),
    to_slogic(92),
    to_slogic(94),
    to_slogic(92),
    to_slogic(99),
    to_slogic(92),
    to_slogic(92),
    to_slogic(81),
    to_slogic(81),
    to_slogic(76),
    to_slogic(81),
    to_slogic(121),
    to_slogic(135),
    to_slogic(151),
    to_slogic(157),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(157),
    to_slogic(144),
    to_slogic(130),
    to_slogic(99),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(89),
    to_slogic(92),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(99),
    to_slogic(89),
    to_slogic(89),
    to_slogic(82),
    to_slogic(176),
    to_slogic(183),
    to_slogic(166),
    to_slogic(146),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(119),
    to_slogic(144),
    to_slogic(83),
    to_slogic(56),
    to_slogic(42),
    to_slogic(50),
    to_slogic(76),
    to_slogic(89),
    to_slogic(56),
    to_slogic(50),
    to_slogic(83),
    to_slogic(65),
    to_slogic(42),
    to_slogic(44),
    to_slogic(97),
    to_slogic(102),
    to_slogic(91),
    to_slogic(102),
    to_slogic(50),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(42),
    to_slogic(68),
    to_slogic(102),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(58),
    to_slogic(87),
    to_slogic(137),
    to_slogic(109),
    to_slogic(185),
    to_slogic(173),
    to_slogic(171),
    to_slogic(182),
    to_slogic(185),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(193),
    to_slogic(118),
    to_slogic(92),
    to_slogic(81),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(96),
    to_slogic(63),
    to_slogic(87),
    to_slogic(63),
    to_slogic(49),
    to_slogic(87),
    to_slogic(75),
    to_slogic(192),
    to_slogic(197),
    to_slogic(193),
    to_slogic(141),
    to_slogic(77),
    to_slogic(102),
    to_slogic(99),
    to_slogic(109),
    to_slogic(118),
    to_slogic(118),
    to_slogic(126),
    to_slogic(134),
    to_slogic(139),
    to_slogic(146),
    to_slogic(151),
    to_slogic(176),
    to_slogic(195),
    to_slogic(213),
    to_slogic(211),
    to_slogic(150),
    to_slogic(82),
    to_slogic(49),
    to_slogic(69),
    to_slogic(49),
    to_slogic(49),
    to_slogic(87),
    to_slogic(96),
    to_slogic(160),
    to_slogic(143),
    to_slogic(92),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(75),
    to_slogic(50),
    to_slogic(126),
    to_slogic(172),
    to_slogic(127),
    to_slogic(87),
    to_slogic(68),
    to_slogic(75),
    to_slogic(63),
    to_slogic(64),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(87),
    to_slogic(132),
    to_slogic(143),
    to_slogic(139),
    to_slogic(139),
    to_slogic(155),
    to_slogic(162),
    to_slogic(158),
    to_slogic(155),
    to_slogic(162),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(157),
    to_slogic(149),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(152),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(132),
    to_slogic(133),
    to_slogic(132),
    to_slogic(133),
    to_slogic(132),
    to_slogic(132),
    to_slogic(100),
    to_slogic(102),
    to_slogic(99),
    to_slogic(96),
    to_slogic(99),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(82),
    to_slogic(81),
    to_slogic(76),
    to_slogic(81),
    to_slogic(116),
    to_slogic(135),
    to_slogic(144),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(157),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(81),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(99),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(63),
    to_slogic(63),
    to_slogic(156),
    to_slogic(109),
    to_slogic(124),
    to_slogic(183),
    to_slogic(177),
    to_slogic(157),
    to_slogic(152),
    to_slogic(128),
    to_slogic(82),
    to_slogic(82),
    to_slogic(49),
    to_slogic(42),
    to_slogic(42),
    to_slogic(76),
    to_slogic(102),
    to_slogic(56),
    to_slogic(44),
    to_slogic(71),
    to_slogic(65),
    to_slogic(71),
    to_slogic(50),
    to_slogic(58),
    to_slogic(97),
    to_slogic(103),
    to_slogic(97),
    to_slogic(115),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(107),
    to_slogic(63),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(36),
    to_slogic(56),
    to_slogic(120),
    to_slogic(101),
    to_slogic(152),
    to_slogic(171),
    to_slogic(155),
    to_slogic(162),
    to_slogic(182),
    to_slogic(191),
    to_slogic(204),
    to_slogic(196),
    to_slogic(193),
    to_slogic(139),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(82),
    to_slogic(63),
    to_slogic(44),
    to_slogic(76),
    to_slogic(109),
    to_slogic(96),
    to_slogic(75),
    to_slogic(83),
    to_slogic(83),
    to_slogic(69),
    to_slogic(126),
    to_slogic(208),
    to_slogic(208),
    to_slogic(197),
    to_slogic(179),
    to_slogic(110),
    to_slogic(99),
    to_slogic(115),
    to_slogic(99),
    to_slogic(115),
    to_slogic(109),
    to_slogic(126),
    to_slogic(126),
    to_slogic(139),
    to_slogic(149),
    to_slogic(162),
    to_slogic(176),
    to_slogic(200),
    to_slogic(214),
    to_slogic(198),
    to_slogic(119),
    to_slogic(96),
    to_slogic(82),
    to_slogic(87),
    to_slogic(83),
    to_slogic(83),
    to_slogic(81),
    to_slogic(81),
    to_slogic(171),
    to_slogic(152),
    to_slogic(102),
    to_slogic(62),
    to_slogic(44),
    to_slogic(33),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(40),
    to_slogic(75),
    to_slogic(46),
    to_slogic(120),
    to_slogic(176),
    to_slogic(126),
    to_slogic(87),
    to_slogic(87),
    to_slogic(83),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(101),
    to_slogic(139),
    to_slogic(139),
    to_slogic(137),
    to_slogic(144),
    to_slogic(155),
    to_slogic(156),
    to_slogic(162),
    to_slogic(150),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(157),
    to_slogic(149),
    to_slogic(152),
    to_slogic(149),
    to_slogic(150),
    to_slogic(155),
    to_slogic(157),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(155),
    to_slogic(152),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(143),
    to_slogic(132),
    to_slogic(126),
    to_slogic(130),
    to_slogic(132),
    to_slogic(132),
    to_slogic(133),
    to_slogic(133),
    to_slogic(158),
    to_slogic(100),
    to_slogic(96),
    to_slogic(99),
    to_slogic(100),
    to_slogic(92),
    to_slogic(102),
    to_slogic(89),
    to_slogic(82),
    to_slogic(89),
    to_slogic(76),
    to_slogic(76),
    to_slogic(89),
    to_slogic(109),
    to_slogic(135),
    to_slogic(151),
    to_slogic(157),
    to_slogic(172),
    to_slogic(176),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(89),
    to_slogic(76),
    to_slogic(82),
    to_slogic(89),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(100),
    to_slogic(116),
    to_slogic(81),
    to_slogic(62),
    to_slogic(56),
    to_slogic(49),
    to_slogic(114),
    to_slogic(141),
    to_slogic(165),
    to_slogic(187),
    to_slogic(213),
    to_slogic(204),
    to_slogic(144),
    to_slogic(63),
    to_slogic(40),
    to_slogic(42),
    to_slogic(42),
    to_slogic(42),
    to_slogic(65),
    to_slogic(83),
    to_slogic(65),
    to_slogic(58),
    to_slogic(56),
    to_slogic(76),
    to_slogic(65),
    to_slogic(65),
    to_slogic(76),
    to_slogic(76),
    to_slogic(115),
    to_slogic(103),
    to_slogic(102),
    to_slogic(120),
    to_slogic(50),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(81),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(42),
    to_slogic(56),
    to_slogic(101),
    to_slogic(109),
    to_slogic(110),
    to_slogic(165),
    to_slogic(156),
    to_slogic(170),
    to_slogic(182),
    to_slogic(196),
    to_slogic(204),
    to_slogic(193),
    to_slogic(193),
    to_slogic(143),
    to_slogic(109),
    to_slogic(117),
    to_slogic(128),
    to_slogic(119),
    to_slogic(126),
    to_slogic(102),
    to_slogic(64),
    to_slogic(56),
    to_slogic(102),
    to_slogic(119),
    to_slogic(96),
    to_slogic(69),
    to_slogic(75),
    to_slogic(118),
    to_slogic(192),
    to_slogic(197),
    to_slogic(211),
    to_slogic(195),
    to_slogic(165),
    to_slogic(134),
    to_slogic(102),
    to_slogic(117),
    to_slogic(115),
    to_slogic(121),
    to_slogic(118),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(146),
    to_slogic(165),
    to_slogic(187),
    to_slogic(211),
    to_slogic(213),
    to_slogic(182),
    to_slogic(110),
    to_slogic(119),
    to_slogic(126),
    to_slogic(87),
    to_slogic(96),
    to_slogic(87),
    to_slogic(87),
    to_slogic(152),
    to_slogic(179),
    to_slogic(149),
    to_slogic(99),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(87),
    to_slogic(49),
    to_slogic(110),
    to_slogic(176),
    to_slogic(133),
    to_slogic(83),
    to_slogic(87),
    to_slogic(83),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(63),
    to_slogic(120),
    to_slogic(143),
    to_slogic(139),
    to_slogic(141),
    to_slogic(152),
    to_slogic(156),
    to_slogic(158),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(157),
    to_slogic(149),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(132),
    to_slogic(133),
    to_slogic(133),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(133),
    to_slogic(143),
    to_slogic(156),
    to_slogic(166),
    to_slogic(171),
    to_slogic(100),
    to_slogic(96),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(89),
    to_slogic(75),
    to_slogic(62),
    to_slogic(81),
    to_slogic(109),
    to_slogic(135),
    to_slogic(144),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(157),
    to_slogic(151),
    to_slogic(121),
    to_slogic(115),
    to_slogic(82),
    to_slogic(82),
    to_slogic(89),
    to_slogic(89),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(97),
    to_slogic(81),
    to_slogic(62),
    to_slogic(49),
    to_slogic(87),
    to_slogic(81),
    to_slogic(113),
    to_slogic(157),
    to_slogic(171),
    to_slogic(165),
    to_slogic(207),
    to_slogic(220),
    to_slogic(166),
    to_slogic(64),
    to_slogic(76),
    to_slogic(42),
    to_slogic(42),
    to_slogic(42),
    to_slogic(65),
    to_slogic(107),
    to_slogic(91),
    to_slogic(71),
    to_slogic(56),
    to_slogic(44),
    to_slogic(83),
    to_slogic(76),
    to_slogic(84),
    to_slogic(84),
    to_slogic(78),
    to_slogic(122),
    to_slogic(91),
    to_slogic(102),
    to_slogic(130),
    to_slogic(65),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(40),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(42),
    to_slogic(68),
    to_slogic(139),
    to_slogic(101),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(182),
    to_slogic(189),
    to_slogic(196),
    to_slogic(196),
    to_slogic(189),
    to_slogic(137),
    to_slogic(116),
    to_slogic(119),
    to_slogic(124),
    to_slogic(126),
    to_slogic(139),
    to_slogic(134),
    to_slogic(128),
    to_slogic(102),
    to_slogic(82),
    to_slogic(102),
    to_slogic(110),
    to_slogic(133),
    to_slogic(128),
    to_slogic(141),
    to_slogic(176),
    to_slogic(191),
    to_slogic(197),
    to_slogic(200),
    to_slogic(187),
    to_slogic(151),
    to_slogic(146),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(118),
    to_slogic(118),
    to_slogic(134),
    to_slogic(126),
    to_slogic(134),
    to_slogic(146),
    to_slogic(165),
    to_slogic(193),
    to_slogic(214),
    to_slogic(214),
    to_slogic(172),
    to_slogic(109),
    to_slogic(102),
    to_slogic(128),
    to_slogic(126),
    to_slogic(113),
    to_slogic(118),
    to_slogic(145),
    to_slogic(179),
    to_slogic(171),
    to_slogic(134),
    to_slogic(99),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(87),
    to_slogic(50),
    to_slogic(101),
    to_slogic(176),
    to_slogic(143),
    to_slogic(83),
    to_slogic(87),
    to_slogic(81),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(83),
    to_slogic(125),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(149),
    to_slogic(162),
    to_slogic(156),
    to_slogic(158),
    to_slogic(150),
    to_slogic(157),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(157),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(151),
    to_slogic(149),
    to_slogic(150),
    to_slogic(152),
    to_slogic(144),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(139),
    to_slogic(143),
    to_slogic(133),
    to_slogic(143),
    to_slogic(132),
    to_slogic(133),
    to_slogic(132),
    to_slogic(144),
    to_slogic(149),
    to_slogic(156),
    to_slogic(166),
    to_slogic(171),
    to_slogic(183),
    to_slogic(183),
    to_slogic(109),
    to_slogic(100),
    to_slogic(96),
    to_slogic(100),
    to_slogic(94),
    to_slogic(99),
    to_slogic(92),
    to_slogic(89),
    to_slogic(89),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(115),
    to_slogic(135),
    to_slogic(152),
    to_slogic(157),
    to_slogic(172),
    to_slogic(173),
    to_slogic(176),
    to_slogic(183),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(172),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(102),
    to_slogic(89),
    to_slogic(81),
    to_slogic(89),
    to_slogic(99),
    to_slogic(99),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(102),
    to_slogic(136),
    to_slogic(70),
    to_slogic(44),
    to_slogic(44),
    to_slogic(69),
    to_slogic(126),
    to_slogic(142),
    to_slogic(161),
    to_slogic(155),
    to_slogic(176),
    to_slogic(176),
    to_slogic(183),
    to_slogic(88),
    to_slogic(56),
    to_slogic(42),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(107),
    to_slogic(115),
    to_slogic(102),
    to_slogic(89),
    to_slogic(36),
    to_slogic(42),
    to_slogic(56),
    to_slogic(78),
    to_slogic(76),
    to_slogic(84),
    to_slogic(78),
    to_slogic(84),
    to_slogic(122),
    to_slogic(103),
    to_slogic(107),
    to_slogic(130),
    to_slogic(95),
    to_slogic(63),
    to_slogic(65),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(40),
    to_slogic(33),
    to_slogic(36),
    to_slogic(49),
    to_slogic(124),
    to_slogic(110),
    to_slogic(141),
    to_slogic(193),
    to_slogic(166),
    to_slogic(171),
    to_slogic(185),
    to_slogic(196),
    to_slogic(204),
    to_slogic(189),
    to_slogic(130),
    to_slogic(109),
    to_slogic(117),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(142),
    to_slogic(109),
    to_slogic(119),
    to_slogic(110),
    to_slogic(118),
    to_slogic(128),
    to_slogic(134),
    to_slogic(151),
    to_slogic(165),
    to_slogic(172),
    to_slogic(169),
    to_slogic(172),
    to_slogic(171),
    to_slogic(161),
    to_slogic(149),
    to_slogic(134),
    to_slogic(124),
    to_slogic(126),
    to_slogic(118),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(149),
    to_slogic(165),
    to_slogic(193),
    to_slogic(214),
    to_slogic(220),
    to_slogic(179),
    to_slogic(152),
    to_slogic(133),
    to_slogic(121),
    to_slogic(149),
    to_slogic(142),
    to_slogic(141),
    to_slogic(161),
    to_slogic(157),
    to_slogic(139),
    to_slogic(99),
    to_slogic(62),
    to_slogic(49),
    to_slogic(76),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(83),
    to_slogic(42),
    to_slogic(101),
    to_slogic(172),
    to_slogic(155),
    to_slogic(87),
    to_slogic(81),
    to_slogic(83),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(68),
    to_slogic(101),
    to_slogic(132),
    to_slogic(139),
    to_slogic(132),
    to_slogic(151),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(162),
    to_slogic(150),
    to_slogic(150),
    to_slogic(155),
    to_slogic(143),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(166),
    to_slogic(165),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(139),
    to_slogic(144),
    to_slogic(143),
    to_slogic(133),
    to_slogic(133),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(149),
    to_slogic(156),
    to_slogic(176),
    to_slogic(171),
    to_slogic(183),
    to_slogic(183),
    to_slogic(183),
    to_slogic(191),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(102),
    to_slogic(92),
    to_slogic(89),
    to_slogic(82),
    to_slogic(81),
    to_slogic(81),
    to_slogic(76),
    to_slogic(76),
    to_slogic(109),
    to_slogic(135),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(130),
    to_slogic(115),
    to_slogic(89),
    to_slogic(81),
    to_slogic(82),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(102),
    to_slogic(115),
    to_slogic(109),
    to_slogic(102),
    to_slogic(143),
    to_slogic(70),
    to_slogic(49),
    to_slogic(96),
    to_slogic(134),
    to_slogic(169),
    to_slogic(141),
    to_slogic(134),
    to_slogic(133),
    to_slogic(149),
    to_slogic(149),
    to_slogic(68),
    to_slogic(63),
    to_slogic(56),
    to_slogic(58),
    to_slogic(65),
    to_slogic(117),
    to_slogic(97),
    to_slogic(71),
    to_slogic(58),
    to_slogic(97),
    to_slogic(56),
    to_slogic(42),
    to_slogic(44),
    to_slogic(63),
    to_slogic(91),
    to_slogic(71),
    to_slogic(91),
    to_slogic(58),
    to_slogic(84),
    to_slogic(117),
    to_slogic(115),
    to_slogic(122),
    to_slogic(115),
    to_slogic(91),
    to_slogic(107),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(42),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(33),
    to_slogic(36),
    to_slogic(83),
    to_slogic(130),
    to_slogic(102),
    to_slogic(170),
    to_slogic(172),
    to_slogic(167),
    to_slogic(182),
    to_slogic(193),
    to_slogic(204),
    to_slogic(193),
    to_slogic(130),
    to_slogic(99),
    to_slogic(118),
    to_slogic(126),
    to_slogic(134),
    to_slogic(142),
    to_slogic(139),
    to_slogic(142),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(142),
    to_slogic(139),
    to_slogic(126),
    to_slogic(117),
    to_slogic(110),
    to_slogic(119),
    to_slogic(127),
    to_slogic(119),
    to_slogic(117),
    to_slogic(117),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(151),
    to_slogic(139),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(142),
    to_slogic(157),
    to_slogic(187),
    to_slogic(214),
    to_slogic(220),
    to_slogic(187),
    to_slogic(165),
    to_slogic(151),
    to_slogic(149),
    to_slogic(146),
    to_slogic(119),
    to_slogic(119),
    to_slogic(119),
    to_slogic(102),
    to_slogic(63),
    to_slogic(63),
    to_slogic(81),
    to_slogic(75),
    to_slogic(89),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(33),
    to_slogic(49),
    to_slogic(63),
    to_slogic(83),
    to_slogic(50),
    to_slogic(96),
    to_slogic(162),
    to_slogic(162),
    to_slogic(102),
    to_slogic(83),
    to_slogic(87),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(83),
    to_slogic(109),
    to_slogic(139),
    to_slogic(139),
    to_slogic(130),
    to_slogic(143),
    to_slogic(156),
    to_slogic(162),
    to_slogic(155),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(151),
    to_slogic(150),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(143),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(152),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(141),
    to_slogic(143),
    to_slogic(132),
    to_slogic(141),
    to_slogic(132),
    to_slogic(133),
    to_slogic(143),
    to_slogic(149),
    to_slogic(166),
    to_slogic(176),
    to_slogic(171),
    to_slogic(183),
    to_slogic(183),
    to_slogic(191),
    to_slogic(183),
    to_slogic(191),
    to_slogic(183),
    to_slogic(102),
    to_slogic(100),
    to_slogic(102),
    to_slogic(96),
    to_slogic(100),
    to_slogic(92),
    to_slogic(92),
    to_slogic(81),
    to_slogic(81),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(115),
    to_slogic(135),
    to_slogic(144),
    to_slogic(157),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(183),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(130),
    to_slogic(115),
    to_slogic(89),
    to_slogic(76),
    to_slogic(89),
    to_slogic(89),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(115),
    to_slogic(115),
    to_slogic(109),
    to_slogic(124),
    to_slogic(120),
    to_slogic(109),
    to_slogic(133),
    to_slogic(128),
    to_slogic(143),
    to_slogic(141),
    to_slogic(110),
    to_slogic(87),
    to_slogic(96),
    to_slogic(87),
    to_slogic(71),
    to_slogic(56),
    to_slogic(42),
    to_slogic(42),
    to_slogic(42),
    to_slogic(83),
    to_slogic(132),
    to_slogic(103),
    to_slogic(109),
    to_slogic(117),
    to_slogic(78),
    to_slogic(56),
    to_slogic(50),
    to_slogic(50),
    to_slogic(84),
    to_slogic(76),
    to_slogic(97),
    to_slogic(65),
    to_slogic(76),
    to_slogic(102),
    to_slogic(109),
    to_slogic(122),
    to_slogic(122),
    to_slogic(130),
    to_slogic(81),
    to_slogic(40),
    to_slogic(50),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(33),
    to_slogic(33),
    to_slogic(56),
    to_slogic(139),
    to_slogic(109),
    to_slogic(134),
    to_slogic(177),
    to_slogic(166),
    to_slogic(171),
    to_slogic(189),
    to_slogic(204),
    to_slogic(196),
    to_slogic(137),
    to_slogic(81),
    to_slogic(100),
    to_slogic(126),
    to_slogic(134),
    to_slogic(142),
    to_slogic(149),
    to_slogic(146),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(134),
    to_slogic(142),
    to_slogic(126),
    to_slogic(126),
    to_slogic(142),
    to_slogic(134),
    to_slogic(142),
    to_slogic(146),
    to_slogic(161),
    to_slogic(151),
    to_slogic(151),
    to_slogic(149),
    to_slogic(133),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(139),
    to_slogic(161),
    to_slogic(183),
    to_slogic(208),
    to_slogic(220),
    to_slogic(193),
    to_slogic(169),
    to_slogic(151),
    to_slogic(149),
    to_slogic(139),
    to_slogic(126),
    to_slogic(127),
    to_slogic(119),
    to_slogic(119),
    to_slogic(92),
    to_slogic(82),
    to_slogic(92),
    to_slogic(89),
    to_slogic(89),
    to_slogic(62),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(75),
    to_slogic(50),
    to_slogic(96),
    to_slogic(165),
    to_slogic(165),
    to_slogic(121),
    to_slogic(75),
    to_slogic(83),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(91),
    to_slogic(134),
    to_slogic(139),
    to_slogic(125),
    to_slogic(139),
    to_slogic(155),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(155),
    to_slogic(143),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(133),
    to_slogic(143),
    to_slogic(156),
    to_slogic(166),
    to_slogic(171),
    to_slogic(183),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(102),
    to_slogic(94),
    to_slogic(102),
    to_slogic(92),
    to_slogic(96),
    to_slogic(92),
    to_slogic(89),
    to_slogic(81),
    to_slogic(89),
    to_slogic(76),
    to_slogic(62),
    to_slogic(76),
    to_slogic(109),
    to_slogic(135),
    to_slogic(144),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(176),
    to_slogic(183),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(178),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(109),
    to_slogic(81),
    to_slogic(76),
    to_slogic(89),
    to_slogic(99),
    to_slogic(89),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(99),
    to_slogic(115),
    to_slogic(102),
    to_slogic(152),
    to_slogic(141),
    to_slogic(169),
    to_slogic(157),
    to_slogic(141),
    to_slogic(109),
    to_slogic(75),
    to_slogic(71),
    to_slogic(75),
    to_slogic(89),
    to_slogic(64),
    to_slogic(42),
    to_slogic(42),
    to_slogic(56),
    to_slogic(50),
    to_slogic(58),
    to_slogic(91),
    to_slogic(140),
    to_slogic(132),
    to_slogic(122),
    to_slogic(107),
    to_slogic(71),
    to_slogic(50),
    to_slogic(42),
    to_slogic(71),
    to_slogic(76),
    to_slogic(84),
    to_slogic(107),
    to_slogic(91),
    to_slogic(76),
    to_slogic(91),
    to_slogic(115),
    to_slogic(130),
    to_slogic(115),
    to_slogic(76),
    to_slogic(63),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(42),
    to_slogic(49),
    to_slogic(40),
    to_slogic(36),
    to_slogic(36),
    to_slogic(96),
    to_slogic(137),
    to_slogic(117),
    to_slogic(167),
    to_slogic(166),
    to_slogic(176),
    to_slogic(185),
    to_slogic(196),
    to_slogic(204),
    to_slogic(144),
    to_slogic(81),
    to_slogic(99),
    to_slogic(118),
    to_slogic(117),
    to_slogic(133),
    to_slogic(134),
    to_slogic(146),
    to_slogic(151),
    to_slogic(149),
    to_slogic(151),
    to_slogic(149),
    to_slogic(149),
    to_slogic(152),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(149),
    to_slogic(146),
    to_slogic(149),
    to_slogic(151),
    to_slogic(161),
    to_slogic(161),
    to_slogic(162),
    to_slogic(161),
    to_slogic(161),
    to_slogic(139),
    to_slogic(128),
    to_slogic(142),
    to_slogic(134),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(151),
    to_slogic(187),
    to_slogic(211),
    to_slogic(220),
    to_slogic(197),
    to_slogic(187),
    to_slogic(169),
    to_slogic(151),
    to_slogic(146),
    to_slogic(142),
    to_slogic(139),
    to_slogic(126),
    to_slogic(126),
    to_slogic(115),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(99),
    to_slogic(70),
    to_slogic(62),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(63),
    to_slogic(75),
    to_slogic(42),
    to_slogic(87),
    to_slogic(162),
    to_slogic(171),
    to_slogic(120),
    to_slogic(64),
    to_slogic(75),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(40),
    to_slogic(49),
    to_slogic(96),
    to_slogic(139),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(152),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(152),
    to_slogic(149),
    to_slogic(155),
    to_slogic(143),
    to_slogic(155),
    to_slogic(143),
    to_slogic(155),
    to_slogic(151),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(139),
    to_slogic(144),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(133),
    to_slogic(144),
    to_slogic(166),
    to_slogic(171),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(183),
    to_slogic(191),
    to_slogic(102),
    to_slogic(102),
    to_slogic(92),
    to_slogic(99),
    to_slogic(82),
    to_slogic(89),
    to_slogic(81),
    to_slogic(81),
    to_slogic(81),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(100),
    to_slogic(130),
    to_slogic(151),
    to_slogic(157),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(115),
    to_slogic(89),
    to_slogic(81),
    to_slogic(81),
    to_slogic(89),
    to_slogic(99),
    to_slogic(99),
    to_slogic(99),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(109),
    to_slogic(126),
    to_slogic(151),
    to_slogic(151),
    to_slogic(117),
    to_slogic(117),
    to_slogic(87),
    to_slogic(64),
    to_slogic(75),
    to_slogic(91),
    to_slogic(71),
    to_slogic(56),
    to_slogic(42),
    to_slogic(65),
    to_slogic(65),
    to_slogic(65),
    to_slogic(78),
    to_slogic(97),
    to_slogic(91),
    to_slogic(89),
    to_slogic(95),
    to_slogic(83),
    to_slogic(42),
    to_slogic(42),
    to_slogic(50),
    to_slogic(58),
    to_slogic(76),
    to_slogic(58),
    to_slogic(97),
    to_slogic(117),
    to_slogic(109),
    to_slogic(109),
    to_slogic(78),
    to_slogic(107),
    to_slogic(81),
    to_slogic(95),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(64),
    to_slogic(143),
    to_slogic(109),
    to_slogic(133),
    to_slogic(171),
    to_slogic(182),
    to_slogic(182),
    to_slogic(193),
    to_slogic(204),
    to_slogic(156),
    to_slogic(76),
    to_slogic(99),
    to_slogic(115),
    to_slogic(115),
    to_slogic(126),
    to_slogic(134),
    to_slogic(142),
    to_slogic(149),
    to_slogic(149),
    to_slogic(151),
    to_slogic(151),
    to_slogic(161),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(149),
    to_slogic(161),
    to_slogic(157),
    to_slogic(161),
    to_slogic(169),
    to_slogic(165),
    to_slogic(169),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(155),
    to_slogic(142),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(157),
    to_slogic(175),
    to_slogic(208),
    to_slogic(220),
    to_slogic(197),
    to_slogic(187),
    to_slogic(169),
    to_slogic(157),
    to_slogic(157),
    to_slogic(149),
    to_slogic(146),
    to_slogic(127),
    to_slogic(128),
    to_slogic(119),
    to_slogic(115),
    to_slogic(119),
    to_slogic(109),
    to_slogic(100),
    to_slogic(76),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(49),
    to_slogic(81),
    to_slogic(158),
    to_slogic(179),
    to_slogic(126),
    to_slogic(63),
    to_slogic(83),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(109),
    to_slogic(139),
    to_slogic(139),
    to_slogic(132),
    to_slogic(144),
    to_slogic(156),
    to_slogic(158),
    to_slogic(155),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(143),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(151),
    to_slogic(143),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(150),
    to_slogic(171),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(102),
    to_slogic(92),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(81),
    to_slogic(82),
    to_slogic(81),
    to_slogic(76),
    to_slogic(62),
    to_slogic(56),
    to_slogic(76),
    to_slogic(100),
    to_slogic(130),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(183),
    to_slogic(178),
    to_slogic(178),
    to_slogic(165),
    to_slogic(151),
    to_slogic(130),
    to_slogic(109),
    to_slogic(89),
    to_slogic(76),
    to_slogic(89),
    to_slogic(99),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(115),
    to_slogic(118),
    to_slogic(119),
    to_slogic(121),
    to_slogic(117),
    to_slogic(117),
    to_slogic(96),
    to_slogic(91),
    to_slogic(109),
    to_slogic(107),
    to_slogic(81),
    to_slogic(50),
    to_slogic(50),
    to_slogic(42),
    to_slogic(76),
    to_slogic(84),
    to_slogic(91),
    to_slogic(109),
    to_slogic(115),
    to_slogic(76),
    to_slogic(65),
    to_slogic(107),
    to_slogic(65),
    to_slogic(40),
    to_slogic(42),
    to_slogic(50),
    to_slogic(76),
    to_slogic(102),
    to_slogic(76),
    to_slogic(58),
    to_slogic(115),
    to_slogic(130),
    to_slogic(103),
    to_slogic(71),
    to_slogic(103),
    to_slogic(145),
    to_slogic(71),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(49),
    to_slogic(118),
    to_slogic(126),
    to_slogic(101),
    to_slogic(162),
    to_slogic(177),
    to_slogic(182),
    to_slogic(189),
    to_slogic(204),
    to_slogic(183),
    to_slogic(76),
    to_slogic(81),
    to_slogic(99),
    to_slogic(115),
    to_slogic(118),
    to_slogic(134),
    to_slogic(142),
    to_slogic(134),
    to_slogic(149),
    to_slogic(149),
    to_slogic(157),
    to_slogic(151),
    to_slogic(172),
    to_slogic(162),
    to_slogic(161),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(169),
    to_slogic(169),
    to_slogic(169),
    to_slogic(165),
    to_slogic(165),
    to_slogic(149),
    to_slogic(139),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(134),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(149),
    to_slogic(187),
    to_slogic(204),
    to_slogic(214),
    to_slogic(211),
    to_slogic(185),
    to_slogic(187),
    to_slogic(165),
    to_slogic(157),
    to_slogic(152),
    to_slogic(149),
    to_slogic(139),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(118),
    to_slogic(102),
    to_slogic(81),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(63),
    to_slogic(63),
    to_slogic(69),
    to_slogic(46),
    to_slogic(81),
    to_slogic(155),
    to_slogic(176),
    to_slogic(133),
    to_slogic(69),
    to_slogic(75),
    to_slogic(44),
    to_slogic(62),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(69),
    to_slogic(118),
    to_slogic(139),
    to_slogic(130),
    to_slogic(139),
    to_slogic(155),
    to_slogic(162),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(152),
    to_slogic(149),
    to_slogic(151),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(143),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(149),
    to_slogic(144),
    to_slogic(139),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(156),
    to_slogic(171),
    to_slogic(183),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(183),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(89),
    to_slogic(89),
    to_slogic(92),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(81),
    to_slogic(76),
    to_slogic(76),
    to_slogic(62),
    to_slogic(56),
    to_slogic(76),
    to_slogic(100),
    to_slogic(130),
    to_slogic(144),
    to_slogic(157),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(115),
    to_slogic(89),
    to_slogic(76),
    to_slogic(81),
    to_slogic(89),
    to_slogic(99),
    to_slogic(99),
    to_slogic(109),
    to_slogic(102),
    to_slogic(115),
    to_slogic(110),
    to_slogic(121),
    to_slogic(122),
    to_slogic(118),
    to_slogic(144),
    to_slogic(157),
    to_slogic(140),
    to_slogic(145),
    to_slogic(130),
    to_slogic(95),
    to_slogic(65),
    to_slogic(63),
    to_slogic(65),
    to_slogic(56),
    to_slogic(97),
    to_slogic(78),
    to_slogic(107),
    to_slogic(115),
    to_slogic(97),
    to_slogic(84),
    to_slogic(107),
    to_slogic(95),
    to_slogic(42),
    to_slogic(42),
    to_slogic(42),
    to_slogic(50),
    to_slogic(65),
    to_slogic(97),
    to_slogic(107),
    to_slogic(84),
    to_slogic(91),
    to_slogic(91),
    to_slogic(109),
    to_slogic(132),
    to_slogic(153),
    to_slogic(102),
    to_slogic(75),
    to_slogic(75),
    to_slogic(69),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(75),
    to_slogic(143),
    to_slogic(101),
    to_slogic(133),
    to_slogic(176),
    to_slogic(182),
    to_slogic(189),
    to_slogic(196),
    to_slogic(189),
    to_slogic(82),
    to_slogic(62),
    to_slogic(81),
    to_slogic(102),
    to_slogic(115),
    to_slogic(124),
    to_slogic(126),
    to_slogic(134),
    to_slogic(139),
    to_slogic(146),
    to_slogic(149),
    to_slogic(151),
    to_slogic(157),
    to_slogic(161),
    to_slogic(165),
    to_slogic(173),
    to_slogic(169),
    to_slogic(172),
    to_slogic(169),
    to_slogic(169),
    to_slogic(169),
    to_slogic(169),
    to_slogic(169),
    to_slogic(169),
    to_slogic(172),
    to_slogic(169),
    to_slogic(165),
    to_slogic(157),
    to_slogic(149),
    to_slogic(144),
    to_slogic(142),
    to_slogic(146),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(118),
    to_slogic(126),
    to_slogic(146),
    to_slogic(175),
    to_slogic(204),
    to_slogic(220),
    to_slogic(211),
    to_slogic(193),
    to_slogic(177),
    to_slogic(169),
    to_slogic(157),
    to_slogic(149),
    to_slogic(146),
    to_slogic(139),
    to_slogic(142),
    to_slogic(134),
    to_slogic(126),
    to_slogic(119),
    to_slogic(118),
    to_slogic(109),
    to_slogic(82),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(75),
    to_slogic(36),
    to_slogic(68),
    to_slogic(157),
    to_slogic(176),
    to_slogic(143),
    to_slogic(69),
    to_slogic(70),
    to_slogic(33),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(91),
    to_slogic(134),
    to_slogic(139),
    to_slogic(137),
    to_slogic(139),
    to_slogic(155),
    to_slogic(156),
    to_slogic(158),
    to_slogic(162),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(144),
    to_slogic(150),
    to_slogic(144),
    to_slogic(150),
    to_slogic(151),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(150),
    to_slogic(171),
    to_slogic(183),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(92),
    to_slogic(96),
    to_slogic(96),
    to_slogic(89),
    to_slogic(82),
    to_slogic(81),
    to_slogic(75),
    to_slogic(76),
    to_slogic(76),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(100),
    to_slogic(135),
    to_slogic(144),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(109),
    to_slogic(89),
    to_slogic(76),
    to_slogic(89),
    to_slogic(89),
    to_slogic(99),
    to_slogic(99),
    to_slogic(103),
    to_slogic(110),
    to_slogic(141),
    to_slogic(144),
    to_slogic(155),
    to_slogic(144),
    to_slogic(160),
    to_slogic(155),
    to_slogic(119),
    to_slogic(83),
    to_slogic(71),
    to_slogic(89),
    to_slogic(63),
    to_slogic(56),
    to_slogic(58),
    to_slogic(65),
    to_slogic(65),
    to_slogic(97),
    to_slogic(84),
    to_slogic(109),
    to_slogic(91),
    to_slogic(107),
    to_slogic(122),
    to_slogic(97),
    to_slogic(56),
    to_slogic(42),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(44),
    to_slogic(63),
    to_slogic(84),
    to_slogic(97),
    to_slogic(117),
    to_slogic(115),
    to_slogic(102),
    to_slogic(102),
    to_slogic(71),
    to_slogic(68),
    to_slogic(126),
    to_slogic(109),
    to_slogic(91),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(42),
    to_slogic(42),
    to_slogic(119),
    to_slogic(128),
    to_slogic(109),
    to_slogic(165),
    to_slogic(182),
    to_slogic(189),
    to_slogic(196),
    to_slogic(207),
    to_slogic(102),
    to_slogic(44),
    to_slogic(76),
    to_slogic(89),
    to_slogic(115),
    to_slogic(118),
    to_slogic(118),
    to_slogic(124),
    to_slogic(134),
    to_slogic(142),
    to_slogic(146),
    to_slogic(146),
    to_slogic(151),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(169),
    to_slogic(177),
    to_slogic(169),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(169),
    to_slogic(172),
    to_slogic(172),
    to_slogic(169),
    to_slogic(172),
    to_slogic(157),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(142),
    to_slogic(126),
    to_slogic(134),
    to_slogic(124),
    to_slogic(134),
    to_slogic(142),
    to_slogic(172),
    to_slogic(193),
    to_slogic(220),
    to_slogic(211),
    to_slogic(195),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(151),
    to_slogic(146),
    to_slogic(139),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(126),
    to_slogic(121),
    to_slogic(109),
    to_slogic(81),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(63),
    to_slogic(64),
    to_slogic(46),
    to_slogic(64),
    to_slogic(157),
    to_slogic(171),
    to_slogic(149),
    to_slogic(69),
    to_slogic(56),
    to_slogic(44),
    to_slogic(62),
    to_slogic(40),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(101),
    to_slogic(139),
    to_slogic(137),
    to_slogic(125),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(149),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(150),
    to_slogic(144),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(141),
    to_slogic(132),
    to_slogic(139),
    to_slogic(132),
    to_slogic(132),
    to_slogic(150),
    to_slogic(166),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(198),
    to_slogic(82),
    to_slogic(89),
    to_slogic(83),
    to_slogic(82),
    to_slogic(81),
    to_slogic(82),
    to_slogic(81),
    to_slogic(76),
    to_slogic(70),
    to_slogic(62),
    to_slogic(56),
    to_slogic(76),
    to_slogic(100),
    to_slogic(130),
    to_slogic(144),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(183),
    to_slogic(173),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(109),
    to_slogic(81),
    to_slogic(76),
    to_slogic(81),
    to_slogic(89),
    to_slogic(92),
    to_slogic(109),
    to_slogic(121),
    to_slogic(134),
    to_slogic(134),
    to_slogic(127),
    to_slogic(133),
    to_slogic(122),
    to_slogic(121),
    to_slogic(96),
    to_slogic(64),
    to_slogic(65),
    to_slogic(83),
    to_slogic(71),
    to_slogic(58),
    to_slogic(58),
    to_slogic(65),
    to_slogic(65),
    to_slogic(84),
    to_slogic(84),
    to_slogic(91),
    to_slogic(109),
    to_slogic(122),
    to_slogic(130),
    to_slogic(107),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(42),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(50),
    to_slogic(71),
    to_slogic(83),
    to_slogic(71),
    to_slogic(102),
    to_slogic(81),
    to_slogic(40),
    to_slogic(42),
    to_slogic(68),
    to_slogic(141),
    to_slogic(125),
    to_slogic(91),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(42),
    to_slogic(83),
    to_slogic(143),
    to_slogic(117),
    to_slogic(125),
    to_slogic(176),
    to_slogic(182),
    to_slogic(193),
    to_slogic(207),
    to_slogic(143),
    to_slogic(44),
    to_slogic(44),
    to_slogic(81),
    to_slogic(100),
    to_slogic(115),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(134),
    to_slogic(139),
    to_slogic(149),
    to_slogic(146),
    to_slogic(149),
    to_slogic(151),
    to_slogic(162),
    to_slogic(165),
    to_slogic(172),
    to_slogic(169),
    to_slogic(177),
    to_slogic(177),
    to_slogic(169),
    to_slogic(176),
    to_slogic(172),
    to_slogic(177),
    to_slogic(172),
    to_slogic(169),
    to_slogic(173),
    to_slogic(161),
    to_slogic(162),
    to_slogic(151),
    to_slogic(146),
    to_slogic(146),
    to_slogic(142),
    to_slogic(139),
    to_slogic(130),
    to_slogic(134),
    to_slogic(126),
    to_slogic(130),
    to_slogic(142),
    to_slogic(165),
    to_slogic(197),
    to_slogic(214),
    to_slogic(214),
    to_slogic(198),
    to_slogic(169),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(146),
    to_slogic(142),
    to_slogic(134),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(118),
    to_slogic(82),
    to_slogic(56),
    to_slogic(44),
    to_slogic(63),
    to_slogic(56),
    to_slogic(69),
    to_slogic(70),
    to_slogic(46),
    to_slogic(64),
    to_slogic(144),
    to_slogic(169),
    to_slogic(158),
    to_slogic(91),
    to_slogic(62),
    to_slogic(33),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(40),
    to_slogic(70),
    to_slogic(118),
    to_slogic(139),
    to_slogic(139),
    to_slogic(137),
    to_slogic(155),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(155),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(151),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(132),
    to_slogic(139),
    to_slogic(132),
    to_slogic(132),
    to_slogic(143),
    to_slogic(166),
    to_slogic(183),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(196),
    to_slogic(191),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(198),
    to_slogic(197),
    to_slogic(198),
    to_slogic(82),
    to_slogic(82),
    to_slogic(81),
    to_slogic(81),
    to_slogic(76),
    to_slogic(75),
    to_slogic(75),
    to_slogic(76),
    to_slogic(70),
    to_slogic(56),
    to_slogic(62),
    to_slogic(63),
    to_slogic(100),
    to_slogic(130),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(130),
    to_slogic(115),
    to_slogic(89),
    to_slogic(76),
    to_slogic(81),
    to_slogic(89),
    to_slogic(99),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(118),
    to_slogic(119),
    to_slogic(133),
    to_slogic(110),
    to_slogic(96),
    to_slogic(91),
    to_slogic(84),
    to_slogic(88),
    to_slogic(83),
    to_slogic(69),
    to_slogic(64),
    to_slogic(56),
    to_slogic(65),
    to_slogic(91),
    to_slogic(97),
    to_slogic(65),
    to_slogic(109),
    to_slogic(130),
    to_slogic(122),
    to_slogic(71),
    to_slogic(83),
    to_slogic(50),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(68),
    to_slogic(71),
    to_slogic(64),
    to_slogic(64),
    to_slogic(40),
    to_slogic(40),
    to_slogic(87),
    to_slogic(125),
    to_slogic(125),
    to_slogic(101),
    to_slogic(75),
    to_slogic(42),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(36),
    to_slogic(49),
    to_slogic(119),
    to_slogic(125),
    to_slogic(119),
    to_slogic(165),
    to_slogic(187),
    to_slogic(189),
    to_slogic(193),
    to_slogic(176),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(81),
    to_slogic(99),
    to_slogic(124),
    to_slogic(118),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(149),
    to_slogic(151),
    to_slogic(165),
    to_slogic(161),
    to_slogic(172),
    to_slogic(172),
    to_slogic(177),
    to_slogic(175),
    to_slogic(187),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(162),
    to_slogic(151),
    to_slogic(149),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(142),
    to_slogic(134),
    to_slogic(134),
    to_slogic(124),
    to_slogic(126),
    to_slogic(142),
    to_slogic(162),
    to_slogic(193),
    to_slogic(220),
    to_slogic(220),
    to_slogic(193),
    to_slogic(172),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(149),
    to_slogic(146),
    to_slogic(134),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(109),
    to_slogic(70),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(75),
    to_slogic(69),
    to_slogic(44),
    to_slogic(50),
    to_slogic(141),
    to_slogic(162),
    to_slogic(144),
    to_slogic(109),
    to_slogic(44),
    to_slogic(33),
    to_slogic(44),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(75),
    to_slogic(124),
    to_slogic(143),
    to_slogic(139),
    to_slogic(139),
    to_slogic(156),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(155),
    to_slogic(155),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(143),
    to_slogic(149),
    to_slogic(151),
    to_slogic(151),
    to_slogic(149),
    to_slogic(144),
    to_slogic(150),
    to_slogic(143),
    to_slogic(144),
    to_slogic(149),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(156),
    to_slogic(183),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(197),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(191),
    to_slogic(197),
    to_slogic(191),
    to_slogic(198),
    to_slogic(197),
    to_slogic(207),
    to_slogic(193),
    to_slogic(207),
    to_slogic(81),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(70),
    to_slogic(63),
    to_slogic(56),
    to_slogic(62),
    to_slogic(100),
    to_slogic(130),
    to_slogic(144),
    to_slogic(157),
    to_slogic(172),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(109),
    to_slogic(89),
    to_slogic(76),
    to_slogic(89),
    to_slogic(92),
    to_slogic(94),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(81),
    to_slogic(82),
    to_slogic(84),
    to_slogic(97),
    to_slogic(91),
    to_slogic(88),
    to_slogic(88),
    to_slogic(69),
    to_slogic(65),
    to_slogic(97),
    to_slogic(107),
    to_slogic(58),
    to_slogic(65),
    to_slogic(122),
    to_slogic(117),
    to_slogic(102),
    to_slogic(65),
    to_slogic(83),
    to_slogic(63),
    to_slogic(42),
    to_slogic(49),
    to_slogic(42),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(75),
    to_slogic(36),
    to_slogic(40),
    to_slogic(83),
    to_slogic(127),
    to_slogic(125),
    to_slogic(144),
    to_slogic(75),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(36),
    to_slogic(75),
    to_slogic(137),
    to_slogic(117),
    to_slogic(134),
    to_slogic(189),
    to_slogic(189),
    to_slogic(193),
    to_slogic(193),
    to_slogic(88),
    to_slogic(40),
    to_slogic(44),
    to_slogic(63),
    to_slogic(82),
    to_slogic(115),
    to_slogic(115),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(142),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(169),
    to_slogic(172),
    to_slogic(176),
    to_slogic(172),
    to_slogic(187),
    to_slogic(169),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(144),
    to_slogic(139),
    to_slogic(134),
    to_slogic(124),
    to_slogic(126),
    to_slogic(134),
    to_slogic(139),
    to_slogic(157),
    to_slogic(195),
    to_slogic(214),
    to_slogic(220),
    to_slogic(200),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(149),
    to_slogic(146),
    to_slogic(142),
    to_slogic(127),
    to_slogic(134),
    to_slogic(126),
    to_slogic(124),
    to_slogic(100),
    to_slogic(76),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(75),
    to_slogic(70),
    to_slogic(33),
    to_slogic(49),
    to_slogic(141),
    to_slogic(162),
    to_slogic(151),
    to_slogic(125),
    to_slogic(44),
    to_slogic(44),
    to_slogic(49),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(96),
    to_slogic(130),
    to_slogic(137),
    to_slogic(139),
    to_slogic(143),
    to_slogic(162),
    to_slogic(162),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(144),
    to_slogic(152),
    to_slogic(155),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(137),
    to_slogic(132),
    to_slogic(119),
    to_slogic(150),
    to_slogic(166),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(191),
    to_slogic(197),
    to_slogic(191),
    to_slogic(196),
    to_slogic(197),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(207),
    to_slogic(193),
    to_slogic(207),
    to_slogic(207),
    to_slogic(82),
    to_slogic(75),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(70),
    to_slogic(70),
    to_slogic(63),
    to_slogic(62),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(97),
    to_slogic(126),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(178),
    to_slogic(172),
    to_slogic(173),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(109),
    to_slogic(81),
    to_slogic(81),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(102),
    to_slogic(100),
    to_slogic(115),
    to_slogic(118),
    to_slogic(103),
    to_slogic(82),
    to_slogic(122),
    to_slogic(130),
    to_slogic(107),
    to_slogic(82),
    to_slogic(102),
    to_slogic(88),
    to_slogic(76),
    to_slogic(102),
    to_slogic(97),
    to_slogic(56),
    to_slogic(44),
    to_slogic(65),
    to_slogic(84),
    to_slogic(132),
    to_slogic(97),
    to_slogic(84),
    to_slogic(63),
    to_slogic(63),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(64),
    to_slogic(40),
    to_slogic(49),
    to_slogic(92),
    to_slogic(110),
    to_slogic(101),
    to_slogic(156),
    to_slogic(125),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(33),
    to_slogic(36),
    to_slogic(40),
    to_slogic(118),
    to_slogic(118),
    to_slogic(117),
    to_slogic(158),
    to_slogic(185),
    to_slogic(193),
    to_slogic(204),
    to_slogic(133),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(81),
    to_slogic(99),
    to_slogic(118),
    to_slogic(124),
    to_slogic(118),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(142),
    to_slogic(146),
    to_slogic(152),
    to_slogic(149),
    to_slogic(157),
    to_slogic(162),
    to_slogic(162),
    to_slogic(165),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(162),
    to_slogic(165),
    to_slogic(151),
    to_slogic(149),
    to_slogic(146),
    to_slogic(142),
    to_slogic(139),
    to_slogic(146),
    to_slogic(134),
    to_slogic(134),
    to_slogic(121),
    to_slogic(126),
    to_slogic(134),
    to_slogic(146),
    to_slogic(157),
    to_slogic(179),
    to_slogic(211),
    to_slogic(220),
    to_slogic(204),
    to_slogic(169),
    to_slogic(165),
    to_slogic(157),
    to_slogic(157),
    to_slogic(149),
    to_slogic(149),
    to_slogic(139),
    to_slogic(134),
    to_slogic(126),
    to_slogic(126),
    to_slogic(124),
    to_slogic(102),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(75),
    to_slogic(63),
    to_slogic(36),
    to_slogic(46),
    to_slogic(141),
    to_slogic(172),
    to_slogic(144),
    to_slogic(144),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(107),
    to_slogic(137),
    to_slogic(139),
    to_slogic(137),
    to_slogic(166),
    to_slogic(167),
    to_slogic(162),
    to_slogic(158),
    to_slogic(155),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(151),
    to_slogic(149),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(139),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(132),
    to_slogic(166),
    to_slogic(183),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(196),
    to_slogic(197),
    to_slogic(197),
    to_slogic(205),
    to_slogic(207),
    to_slogic(193),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(193),
    to_slogic(76),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(69),
    to_slogic(70),
    to_slogic(70),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(97),
    to_slogic(134),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(172),
    to_slogic(165),
    to_slogic(143),
    to_slogic(135),
    to_slogic(115),
    to_slogic(81),
    to_slogic(76),
    to_slogic(82),
    to_slogic(103),
    to_slogic(110),
    to_slogic(99),
    to_slogic(100),
    to_slogic(118),
    to_slogic(102),
    to_slogic(117),
    to_slogic(122),
    to_slogic(138),
    to_slogic(126),
    to_slogic(89),
    to_slogic(82),
    to_slogic(102),
    to_slogic(113),
    to_slogic(71),
    to_slogic(115),
    to_slogic(84),
    to_slogic(58),
    to_slogic(76),
    to_slogic(76),
    to_slogic(58),
    to_slogic(76),
    to_slogic(130),
    to_slogic(97),
    to_slogic(107),
    to_slogic(50),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(89),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(87),
    to_slogic(121),
    to_slogic(96),
    to_slogic(118),
    to_slogic(150),
    to_slogic(119),
    to_slogic(49),
    to_slogic(36),
    to_slogic(40),
    to_slogic(40),
    to_slogic(64),
    to_slogic(137),
    to_slogic(109),
    to_slogic(127),
    to_slogic(191),
    to_slogic(193),
    to_slogic(205),
    to_slogic(176),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(81),
    to_slogic(102),
    to_slogic(115),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(151),
    to_slogic(149),
    to_slogic(157),
    to_slogic(162),
    to_slogic(172),
    to_slogic(169),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(157),
    to_slogic(165),
    to_slogic(146),
    to_slogic(144),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(134),
    to_slogic(142),
    to_slogic(149),
    to_slogic(172),
    to_slogic(211),
    to_slogic(220),
    to_slogic(211),
    to_slogic(165),
    to_slogic(162),
    to_slogic(157),
    to_slogic(151),
    to_slogic(146),
    to_slogic(149),
    to_slogic(133),
    to_slogic(142),
    to_slogic(128),
    to_slogic(124),
    to_slogic(118),
    to_slogic(89),
    to_slogic(62),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(82),
    to_slogic(62),
    to_slogic(36),
    to_slogic(36),
    to_slogic(134),
    to_slogic(162),
    to_slogic(144),
    to_slogic(144),
    to_slogic(63),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(75),
    to_slogic(124),
    to_slogic(137),
    to_slogic(137),
    to_slogic(143),
    to_slogic(162),
    to_slogic(166),
    to_slogic(158),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(150),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(139),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(150),
    to_slogic(178),
    to_slogic(191),
    to_slogic(196),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(198),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(193),
    to_slogic(207),
    to_slogic(82),
    to_slogic(75),
    to_slogic(76),
    to_slogic(69),
    to_slogic(75),
    to_slogic(75),
    to_slogic(70),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(100),
    to_slogic(130),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(176),
    to_slogic(172),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(115),
    to_slogic(81),
    to_slogic(76),
    to_slogic(77),
    to_slogic(109),
    to_slogic(117),
    to_slogic(92),
    to_slogic(103),
    to_slogic(117),
    to_slogic(141),
    to_slogic(160),
    to_slogic(141),
    to_slogic(68),
    to_slogic(56),
    to_slogic(63),
    to_slogic(103),
    to_slogic(143),
    to_slogic(84),
    to_slogic(107),
    to_slogic(89),
    to_slogic(50),
    to_slogic(58),
    to_slogic(102),
    to_slogic(78),
    to_slogic(58),
    to_slogic(109),
    to_slogic(132),
    to_slogic(109),
    to_slogic(120),
    to_slogic(71),
    to_slogic(50),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(42),
    to_slogic(49),
    to_slogic(75),
    to_slogic(70),
    to_slogic(64),
    to_slogic(49),
    to_slogic(69),
    to_slogic(96),
    to_slogic(149),
    to_slogic(128),
    to_slogic(70),
    to_slogic(107),
    to_slogic(158),
    to_slogic(83),
    to_slogic(33),
    to_slogic(33),
    to_slogic(36),
    to_slogic(102),
    to_slogic(124),
    to_slogic(117),
    to_slogic(149),
    to_slogic(204),
    to_slogic(204),
    to_slogic(207),
    to_slogic(102),
    to_slogic(40),
    to_slogic(36),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(81),
    to_slogic(99),
    to_slogic(99),
    to_slogic(118),
    to_slogic(124),
    to_slogic(130),
    to_slogic(126),
    to_slogic(134),
    to_slogic(139),
    to_slogic(142),
    to_slogic(146),
    to_slogic(146),
    to_slogic(151),
    to_slogic(157),
    to_slogic(161),
    to_slogic(165),
    to_slogic(161),
    to_slogic(173),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(152),
    to_slogic(149),
    to_slogic(144),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(124),
    to_slogic(118),
    to_slogic(121),
    to_slogic(126),
    to_slogic(134),
    to_slogic(151),
    to_slogic(175),
    to_slogic(211),
    to_slogic(220),
    to_slogic(211),
    to_slogic(169),
    to_slogic(165),
    to_slogic(157),
    to_slogic(151),
    to_slogic(146),
    to_slogic(142),
    to_slogic(139),
    to_slogic(134),
    to_slogic(134),
    to_slogic(126),
    to_slogic(121),
    to_slogic(82),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(75),
    to_slogic(70),
    to_slogic(33),
    to_slogic(46),
    to_slogic(109),
    to_slogic(169),
    to_slogic(141),
    to_slogic(141),
    to_slogic(83),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(83),
    to_slogic(137),
    to_slogic(137),
    to_slogic(137),
    to_slogic(151),
    to_slogic(158),
    to_slogic(162),
    to_slogic(156),
    to_slogic(150),
    to_slogic(158),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(143),
    to_slogic(149),
    to_slogic(151),
    to_slogic(143),
    to_slogic(150),
    to_slogic(144),
    to_slogic(151),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(132),
    to_slogic(144),
    to_slogic(139),
    to_slogic(130),
    to_slogic(130),
    to_slogic(143),
    to_slogic(166),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(193),
    to_slogic(207),
    to_slogic(207),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(70),
    to_slogic(69),
    to_slogic(62),
    to_slogic(56),
    to_slogic(44),
    to_slogic(62),
    to_slogic(97),
    to_slogic(130),
    to_slogic(144),
    to_slogic(151),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(143),
    to_slogic(130),
    to_slogic(109),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(110),
    to_slogic(133),
    to_slogic(103),
    to_slogic(133),
    to_slogic(148),
    to_slogic(133),
    to_slogic(121),
    to_slogic(117),
    to_slogic(50),
    to_slogic(63),
    to_slogic(96),
    to_slogic(126),
    to_slogic(113),
    to_slogic(102),
    to_slogic(81),
    to_slogic(58),
    to_slogic(58),
    to_slogic(78),
    to_slogic(97),
    to_slogic(109),
    to_slogic(65),
    to_slogic(132),
    to_slogic(117),
    to_slogic(122),
    to_slogic(97),
    to_slogic(97),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(82),
    to_slogic(101),
    to_slogic(82),
    to_slogic(63),
    to_slogic(69),
    to_slogic(88),
    to_slogic(121),
    to_slogic(176),
    to_slogic(165),
    to_slogic(75),
    to_slogic(69),
    to_slogic(118),
    to_slogic(75),
    to_slogic(33),
    to_slogic(33),
    to_slogic(56),
    to_slogic(139),
    to_slogic(117),
    to_slogic(119),
    to_slogic(176),
    to_slogic(204),
    to_slogic(204),
    to_slogic(143),
    to_slogic(40),
    to_slogic(33),
    to_slogic(33),
    to_slogic(64),
    to_slogic(70),
    to_slogic(56),
    to_slogic(76),
    to_slogic(99),
    to_slogic(115),
    to_slogic(121),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(162),
    to_slogic(157),
    to_slogic(162),
    to_slogic(157),
    to_slogic(146),
    to_slogic(139),
    to_slogic(134),
    to_slogic(130),
    to_slogic(134),
    to_slogic(134),
    to_slogic(126),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(134),
    to_slogic(149),
    to_slogic(169),
    to_slogic(193),
    to_slogic(220),
    to_slogic(220),
    to_slogic(179),
    to_slogic(157),
    to_slogic(157),
    to_slogic(149),
    to_slogic(146),
    to_slogic(146),
    to_slogic(142),
    to_slogic(134),
    to_slogic(126),
    to_slogic(124),
    to_slogic(102),
    to_slogic(81),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(64),
    to_slogic(75),
    to_slogic(70),
    to_slogic(36),
    to_slogic(44),
    to_slogic(101),
    to_slogic(162),
    to_slogic(143),
    to_slogic(149),
    to_slogic(96),
    to_slogic(33),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(107),
    to_slogic(137),
    to_slogic(137),
    to_slogic(139),
    to_slogic(150),
    to_slogic(162),
    to_slogic(156),
    to_slogic(158),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(143),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(139),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(158),
    to_slogic(183),
    to_slogic(191),
    to_slogic(197),
    to_slogic(196),
    to_slogic(196),
    to_slogic(191),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(193),
    to_slogic(207),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(77),
    to_slogic(75),
    to_slogic(70),
    to_slogic(63),
    to_slogic(62),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(97),
    to_slogic(130),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(176),
    to_slogic(172),
    to_slogic(157),
    to_slogic(151),
    to_slogic(135),
    to_slogic(109),
    to_slogic(81),
    to_slogic(62),
    to_slogic(76),
    to_slogic(92),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(110),
    to_slogic(113),
    to_slogic(128),
    to_slogic(110),
    to_slogic(63),
    to_slogic(81),
    to_slogic(122),
    to_slogic(107),
    to_slogic(83),
    to_slogic(89),
    to_slogic(89),
    to_slogic(76),
    to_slogic(65),
    to_slogic(97),
    to_slogic(91),
    to_slogic(109),
    to_slogic(78),
    to_slogic(130),
    to_slogic(109),
    to_slogic(145),
    to_slogic(89),
    to_slogic(115),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(42),
    to_slogic(33),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(70),
    to_slogic(107),
    to_slogic(82),
    to_slogic(63),
    to_slogic(81),
    to_slogic(110),
    to_slogic(119),
    to_slogic(167),
    to_slogic(171),
    to_slogic(91),
    to_slogic(49),
    to_slogic(88),
    to_slogic(49),
    to_slogic(33),
    to_slogic(33),
    to_slogic(91),
    to_slogic(136),
    to_slogic(119),
    to_slogic(141),
    to_slogic(196),
    to_slogic(196),
    to_slogic(171),
    to_slogic(56),
    to_slogic(33),
    to_slogic(33),
    to_slogic(36),
    to_slogic(64),
    to_slogic(76),
    to_slogic(62),
    to_slogic(76),
    to_slogic(97),
    to_slogic(99),
    to_slogic(118),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(157),
    to_slogic(165),
    to_slogic(151),
    to_slogic(144),
    to_slogic(139),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(118),
    to_slogic(124),
    to_slogic(134),
    to_slogic(149),
    to_slogic(165),
    to_slogic(187),
    to_slogic(220),
    to_slogic(220),
    to_slogic(187),
    to_slogic(155),
    to_slogic(151),
    to_slogic(151),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(127),
    to_slogic(134),
    to_slogic(121),
    to_slogic(100),
    to_slogic(63),
    to_slogic(46),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(64),
    to_slogic(70),
    to_slogic(70),
    to_slogic(33),
    to_slogic(44),
    to_slogic(87),
    to_slogic(165),
    to_slogic(151),
    to_slogic(149),
    to_slogic(102),
    to_slogic(33),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(63),
    to_slogic(118),
    to_slogic(139),
    to_slogic(137),
    to_slogic(137),
    to_slogic(158),
    to_slogic(156),
    to_slogic(158),
    to_slogic(162),
    to_slogic(157),
    to_slogic(152),
    to_slogic(158),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(144),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(132),
    to_slogic(144),
    to_slogic(139),
    to_slogic(132),
    to_slogic(132),
    to_slogic(143),
    to_slogic(166),
    to_slogic(191),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(191),
    to_slogic(197),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(82),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(69),
    to_slogic(75),
    to_slogic(70),
    to_slogic(70),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(97),
    to_slogic(130),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(161),
    to_slogic(151),
    to_slogic(135),
    to_slogic(109),
    to_slogic(81),
    to_slogic(76),
    to_slogic(76),
    to_slogic(81),
    to_slogic(96),
    to_slogic(110),
    to_slogic(121),
    to_slogic(122),
    to_slogic(122),
    to_slogic(133),
    to_slogic(121),
    to_slogic(63),
    to_slogic(69),
    to_slogic(102),
    to_slogic(96),
    to_slogic(91),
    to_slogic(91),
    to_slogic(78),
    to_slogic(65),
    to_slogic(91),
    to_slogic(78),
    to_slogic(117),
    to_slogic(97),
    to_slogic(78),
    to_slogic(109),
    to_slogic(109),
    to_slogic(145),
    to_slogic(76),
    to_slogic(102),
    to_slogic(50),
    to_slogic(40),
    to_slogic(42),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(63),
    to_slogic(81),
    to_slogic(83),
    to_slogic(82),
    to_slogic(91),
    to_slogic(139),
    to_slogic(107),
    to_slogic(81),
    to_slogic(88),
    to_slogic(124),
    to_slogic(82),
    to_slogic(33),
    to_slogic(56),
    to_slogic(33),
    to_slogic(33),
    to_slogic(49),
    to_slogic(124),
    to_slogic(117),
    to_slogic(119),
    to_slogic(177),
    to_slogic(207),
    to_slogic(193),
    to_slogic(82),
    to_slogic(33),
    to_slogic(40),
    to_slogic(44),
    to_slogic(33),
    to_slogic(75),
    to_slogic(81),
    to_slogic(62),
    to_slogic(76),
    to_slogic(97),
    to_slogic(115),
    to_slogic(121),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(142),
    to_slogic(146),
    to_slogic(149),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(162),
    to_slogic(162),
    to_slogic(151),
    to_slogic(162),
    to_slogic(157),
    to_slogic(146),
    to_slogic(144),
    to_slogic(134),
    to_slogic(130),
    to_slogic(124),
    to_slogic(126),
    to_slogic(139),
    to_slogic(126),
    to_slogic(118),
    to_slogic(124),
    to_slogic(118),
    to_slogic(134),
    to_slogic(144),
    to_slogic(161),
    to_slogic(179),
    to_slogic(220),
    to_slogic(226),
    to_slogic(195),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(149),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(126),
    to_slogic(117),
    to_slogic(92),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(64),
    to_slogic(75),
    to_slogic(70),
    to_slogic(33),
    to_slogic(36),
    to_slogic(83),
    to_slogic(155),
    to_slogic(149),
    to_slogic(155),
    to_slogic(109),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(83),
    to_slogic(124),
    to_slogic(137),
    to_slogic(144),
    to_slogic(143),
    to_slogic(162),
    to_slogic(156),
    to_slogic(158),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(149),
    to_slogic(143),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(158),
    to_slogic(183),
    to_slogic(196),
    to_slogic(197),
    to_slogic(197),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(191),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(82),
    to_slogic(75),
    to_slogic(81),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(70),
    to_slogic(63),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(89),
    to_slogic(121),
    to_slogic(144),
    to_slogic(157),
    to_slogic(162),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(165),
    to_slogic(143),
    to_slogic(135),
    to_slogic(115),
    to_slogic(81),
    to_slogic(76),
    to_slogic(76),
    to_slogic(82),
    to_slogic(103),
    to_slogic(117),
    to_slogic(121),
    to_slogic(110),
    to_slogic(121),
    to_slogic(128),
    to_slogic(88),
    to_slogic(63),
    to_slogic(88),
    to_slogic(82),
    to_slogic(84),
    to_slogic(107),
    to_slogic(84),
    to_slogic(76),
    to_slogic(91),
    to_slogic(76),
    to_slogic(78),
    to_slogic(120),
    to_slogic(58),
    to_slogic(78),
    to_slogic(103),
    to_slogic(102),
    to_slogic(155),
    to_slogic(84),
    to_slogic(83),
    to_slogic(71),
    to_slogic(40),
    to_slogic(49),
    to_slogic(42),
    to_slogic(56),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(81),
    to_slogic(63),
    to_slogic(83),
    to_slogic(125),
    to_slogic(130),
    to_slogic(96),
    to_slogic(77),
    to_slogic(102),
    to_slogic(83),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(33),
    to_slogic(68),
    to_slogic(96),
    to_slogic(118),
    to_slogic(117),
    to_slogic(132),
    to_slogic(189),
    to_slogic(156),
    to_slogic(130),
    to_slogic(49),
    to_slogic(33),
    to_slogic(33),
    to_slogic(44),
    to_slogic(33),
    to_slogic(82),
    to_slogic(83),
    to_slogic(62),
    to_slogic(76),
    to_slogic(97),
    to_slogic(99),
    to_slogic(115),
    to_slogic(118),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(152),
    to_slogic(149),
    to_slogic(152),
    to_slogic(149),
    to_slogic(157),
    to_slogic(161),
    to_slogic(165),
    to_slogic(151),
    to_slogic(162),
    to_slogic(151),
    to_slogic(149),
    to_slogic(146),
    to_slogic(144),
    to_slogic(126),
    to_slogic(115),
    to_slogic(118),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(134),
    to_slogic(142),
    to_slogic(162),
    to_slogic(176),
    to_slogic(214),
    to_slogic(226),
    to_slogic(200),
    to_slogic(152),
    to_slogic(146),
    to_slogic(151),
    to_slogic(146),
    to_slogic(146),
    to_slogic(134),
    to_slogic(128),
    to_slogic(126),
    to_slogic(117),
    to_slogic(75),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(75),
    to_slogic(64),
    to_slogic(62),
    to_slogic(44),
    to_slogic(33),
    to_slogic(77),
    to_slogic(143),
    to_slogic(157),
    to_slogic(149),
    to_slogic(126),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(96),
    to_slogic(137),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(152),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(151),
    to_slogic(150),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(139),
    to_slogic(132),
    to_slogic(137),
    to_slogic(132),
    to_slogic(144),
    to_slogic(166),
    to_slogic(191),
    to_slogic(197),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(205),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(89),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(75),
    to_slogic(70),
    to_slogic(70),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(33),
    to_slogic(56),
    to_slogic(89),
    to_slogic(130),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(115),
    to_slogic(81),
    to_slogic(69),
    to_slogic(82),
    to_slogic(110),
    to_slogic(133),
    to_slogic(117),
    to_slogic(102),
    to_slogic(110),
    to_slogic(110),
    to_slogic(110),
    to_slogic(81),
    to_slogic(69),
    to_slogic(84),
    to_slogic(82),
    to_slogic(97),
    to_slogic(115),
    to_slogic(75),
    to_slogic(84),
    to_slogic(76),
    to_slogic(58),
    to_slogic(115),
    to_slogic(91),
    to_slogic(44),
    to_slogic(97),
    to_slogic(109),
    to_slogic(91),
    to_slogic(145),
    to_slogic(103),
    to_slogic(68),
    to_slogic(97),
    to_slogic(42),
    to_slogic(50),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(63),
    to_slogic(81),
    to_slogic(130),
    to_slogic(101),
    to_slogic(92),
    to_slogic(118),
    to_slogic(124),
    to_slogic(83),
    to_slogic(64),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(36),
    to_slogic(49),
    to_slogic(143),
    to_slogic(151),
    to_slogic(130),
    to_slogic(114),
    to_slogic(120),
    to_slogic(156),
    to_slogic(167),
    to_slogic(118),
    to_slogic(49),
    to_slogic(44),
    to_slogic(33),
    to_slogic(33),
    to_slogic(49),
    to_slogic(75),
    to_slogic(94),
    to_slogic(76),
    to_slogic(76),
    to_slogic(89),
    to_slogic(115),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(146),
    to_slogic(139),
    to_slogic(118),
    to_slogic(115),
    to_slogic(118),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(124),
    to_slogic(126),
    to_slogic(139),
    to_slogic(157),
    to_slogic(179),
    to_slogic(211),
    to_slogic(226),
    to_slogic(200),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(134),
    to_slogic(126),
    to_slogic(124),
    to_slogic(109),
    to_slogic(56),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(64),
    to_slogic(75),
    to_slogic(62),
    to_slogic(44),
    to_slogic(33),
    to_slogic(56),
    to_slogic(144),
    to_slogic(162),
    to_slogic(155),
    to_slogic(139),
    to_slogic(64),
    to_slogic(49),
    to_slogic(36),
    to_slogic(56),
    to_slogic(109),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(149),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(155),
    to_slogic(143),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(150),
    to_slogic(143),
    to_slogic(149),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(137),
    to_slogic(125),
    to_slogic(132),
    to_slogic(158),
    to_slogic(183),
    to_slogic(191),
    to_slogic(197),
    to_slogic(196),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(82),
    to_slogic(82),
    to_slogic(75),
    to_slogic(81),
    to_slogic(75),
    to_slogic(76),
    to_slogic(70),
    to_slogic(70),
    to_slogic(62),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(100),
    to_slogic(121),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(176),
    to_slogic(172),
    to_slogic(165),
    to_slogic(151),
    to_slogic(130),
    to_slogic(115),
    to_slogic(82),
    to_slogic(103),
    to_slogic(121),
    to_slogic(127),
    to_slogic(109),
    to_slogic(102),
    to_slogic(102),
    to_slogic(110),
    to_slogic(124),
    to_slogic(110),
    to_slogic(75),
    to_slogic(69),
    to_slogic(82),
    to_slogic(91),
    to_slogic(122),
    to_slogic(102),
    to_slogic(76),
    to_slogic(65),
    to_slogic(58),
    to_slogic(76),
    to_slogic(122),
    to_slogic(76),
    to_slogic(44),
    to_slogic(84),
    to_slogic(109),
    to_slogic(78),
    to_slogic(143),
    to_slogic(115),
    to_slogic(56),
    to_slogic(122),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(33),
    to_slogic(49),
    to_slogic(68),
    to_slogic(75),
    to_slogic(56),
    to_slogic(40),
    to_slogic(69),
    to_slogic(110),
    to_slogic(83),
    to_slogic(33),
    to_slogic(33),
    to_slogic(33),
    to_slogic(40),
    to_slogic(33),
    to_slogic(102),
    to_slogic(158),
    to_slogic(167),
    to_slogic(167),
    to_slogic(165),
    to_slogic(167),
    to_slogic(176),
    to_slogic(143),
    to_slogic(64),
    to_slogic(33),
    to_slogic(33),
    to_slogic(49),
    to_slogic(44),
    to_slogic(33),
    to_slogic(82),
    to_slogic(96),
    to_slogic(62),
    to_slogic(76),
    to_slogic(97),
    to_slogic(115),
    to_slogic(115),
    to_slogic(118),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(152),
    to_slogic(149),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(126),
    to_slogic(115),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(130),
    to_slogic(139),
    to_slogic(134),
    to_slogic(124),
    to_slogic(118),
    to_slogic(134),
    to_slogic(152),
    to_slogic(177),
    to_slogic(200),
    to_slogic(211),
    to_slogic(187),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(142),
    to_slogic(128),
    to_slogic(128),
    to_slogic(117),
    to_slogic(82),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(64),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(133),
    to_slogic(162),
    to_slogic(149),
    to_slogic(133),
    to_slogic(83),
    to_slogic(40),
    to_slogic(40),
    to_slogic(63),
    to_slogic(125),
    to_slogic(152),
    to_slogic(137),
    to_slogic(143),
    to_slogic(157),
    to_slogic(162),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(158),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(152),
    to_slogic(149),
    to_slogic(150),
    to_slogic(151),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(132),
    to_slogic(139),
    to_slogic(132),
    to_slogic(132),
    to_slogic(139),
    to_slogic(166),
    to_slogic(191),
    to_slogic(197),
    to_slogic(196),
    to_slogic(191),
    to_slogic(196),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(205),
    to_slogic(193),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(76),
    to_slogic(62),
    to_slogic(62),
    to_slogic(62),
    to_slogic(44),
    to_slogic(62),
    to_slogic(100),
    to_slogic(134),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(117),
    to_slogic(103),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(102),
    to_slogic(99),
    to_slogic(110),
    to_slogic(121),
    to_slogic(110),
    to_slogic(81),
    to_slogic(63),
    to_slogic(88),
    to_slogic(91),
    to_slogic(115),
    to_slogic(102),
    to_slogic(76),
    to_slogic(50),
    to_slogic(58),
    to_slogic(130),
    to_slogic(107),
    to_slogic(65),
    to_slogic(58),
    to_slogic(71),
    to_slogic(117),
    to_slogic(86),
    to_slogic(130),
    to_slogic(153),
    to_slogic(65),
    to_slogic(127),
    to_slogic(71),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(36),
    to_slogic(40),
    to_slogic(63),
    to_slogic(56),
    to_slogic(50),
    to_slogic(56),
    to_slogic(113),
    to_slogic(87),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(36),
    to_slogic(36),
    to_slogic(149),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(182),
    to_slogic(176),
    to_slogic(143),
    to_slogic(75),
    to_slogic(33),
    to_slogic(33),
    to_slogic(33),
    to_slogic(49),
    to_slogic(44),
    to_slogic(36),
    to_slogic(82),
    to_slogic(96),
    to_slogic(76),
    to_slogic(76),
    to_slogic(97),
    to_slogic(109),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(152),
    to_slogic(149),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(146),
    to_slogic(139),
    to_slogic(134),
    to_slogic(115),
    to_slogic(130),
    to_slogic(130),
    to_slogic(97),
    to_slogic(76),
    to_slogic(89),
    to_slogic(115),
    to_slogic(115),
    to_slogic(115),
    to_slogic(124),
    to_slogic(139),
    to_slogic(165),
    to_slogic(193),
    to_slogic(195),
    to_slogic(162),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(146),
    to_slogic(139),
    to_slogic(134),
    to_slogic(124),
    to_slogic(109),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(42),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(70),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(33),
    to_slogic(44),
    to_slogic(120),
    to_slogic(162),
    to_slogic(157),
    to_slogic(132),
    to_slogic(83),
    to_slogic(44),
    to_slogic(40),
    to_slogic(75),
    to_slogic(137),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(162),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(143),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(139),
    to_slogic(139),
    to_slogic(125),
    to_slogic(150),
    to_slogic(166),
    to_slogic(191),
    to_slogic(197),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(191),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(82),
    to_slogic(75),
    to_slogic(81),
    to_slogic(76),
    to_slogic(75),
    to_slogic(81),
    to_slogic(70),
    to_slogic(62),
    to_slogic(62),
    to_slogic(62),
    to_slogic(56),
    to_slogic(76),
    to_slogic(115),
    to_slogic(133),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(152),
    to_slogic(135),
    to_slogic(126),
    to_slogic(82),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(99),
    to_slogic(102),
    to_slogic(110),
    to_slogic(110),
    to_slogic(87),
    to_slogic(81),
    to_slogic(69),
    to_slogic(96),
    to_slogic(91),
    to_slogic(134),
    to_slogic(96),
    to_slogic(71),
    to_slogic(42),
    to_slogic(76),
    to_slogic(130),
    to_slogic(76),
    to_slogic(83),
    to_slogic(76),
    to_slogic(71),
    to_slogic(109),
    to_slogic(86),
    to_slogic(122),
    to_slogic(155),
    to_slogic(84),
    to_slogic(102),
    to_slogic(89),
    to_slogic(40),
    to_slogic(42),
    to_slogic(82),
    to_slogic(64),
    to_slogic(56),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(42),
    to_slogic(76),
    to_slogic(81),
    to_slogic(153),
    to_slogic(69),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(63),
    to_slogic(158),
    to_slogic(167),
    to_slogic(189),
    to_slogic(189),
    to_slogic(193),
    to_slogic(167),
    to_slogic(64),
    to_slogic(33),
    to_slogic(33),
    to_slogic(33),
    to_slogic(40),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(75),
    to_slogic(109),
    to_slogic(76),
    to_slogic(97),
    to_slogic(97),
    to_slogic(115),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(149),
    to_slogic(146),
    to_slogic(146),
    to_slogic(134),
    to_slogic(118),
    to_slogic(130),
    to_slogic(130),
    to_slogic(97),
    to_slogic(77),
    to_slogic(97),
    to_slogic(99),
    to_slogic(97),
    to_slogic(99),
    to_slogic(115),
    to_slogic(124),
    to_slogic(151),
    to_slogic(187),
    to_slogic(187),
    to_slogic(165),
    to_slogic(151),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(134),
    to_slogic(134),
    to_slogic(124),
    to_slogic(82),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(70),
    to_slogic(70),
    to_slogic(75),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(36),
    to_slogic(101),
    to_slogic(165),
    to_slogic(149),
    to_slogic(141),
    to_slogic(91),
    to_slogic(40),
    to_slogic(56),
    to_slogic(96),
    to_slogic(137),
    to_slogic(152),
    to_slogic(144),
    to_slogic(150),
    to_slogic(162),
    to_slogic(150),
    to_slogic(158),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(151),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(144),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(158),
    to_slogic(183),
    to_slogic(191),
    to_slogic(197),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(75),
    to_slogic(82),
    to_slogic(81),
    to_slogic(75),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(62),
    to_slogic(70),
    to_slogic(70),
    to_slogic(62),
    to_slogic(82),
    to_slogic(117),
    to_slogic(139),
    to_slogic(152),
    to_slogic(157),
    to_slogic(162),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(135),
    to_slogic(115),
    to_slogic(82),
    to_slogic(76),
    to_slogic(81),
    to_slogic(92),
    to_slogic(99),
    to_slogic(100),
    to_slogic(102),
    to_slogic(110),
    to_slogic(117),
    to_slogic(103),
    to_slogic(88),
    to_slogic(69),
    to_slogic(91),
    to_slogic(82),
    to_slogic(88),
    to_slogic(71),
    to_slogic(58),
    to_slogic(50),
    to_slogic(122),
    to_slogic(107),
    to_slogic(65),
    to_slogic(91),
    to_slogic(78),
    to_slogic(58),
    to_slogic(122),
    to_slogic(97),
    to_slogic(109),
    to_slogic(143),
    to_slogic(109),
    to_slogic(95),
    to_slogic(120),
    to_slogic(33),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(124),
    to_slogic(82),
    to_slogic(40),
    to_slogic(36),
    to_slogic(36),
    to_slogic(56),
    to_slogic(113),
    to_slogic(87),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(69),
    to_slogic(101),
    to_slogic(139),
    to_slogic(150),
    to_slogic(162),
    to_slogic(171),
    to_slogic(171),
    to_slogic(102),
    to_slogic(33),
    to_slogic(33),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(46),
    to_slogic(82),
    to_slogic(109),
    to_slogic(76),
    to_slogic(97),
    to_slogic(97),
    to_slogic(115),
    to_slogic(115),
    to_slogic(118),
    to_slogic(124),
    to_slogic(118),
    to_slogic(124),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(142),
    to_slogic(144),
    to_slogic(142),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(151),
    to_slogic(149),
    to_slogic(152),
    to_slogic(161),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(146),
    to_slogic(146),
    to_slogic(126),
    to_slogic(124),
    to_slogic(118),
    to_slogic(124),
    to_slogic(130),
    to_slogic(126),
    to_slogic(124),
    to_slogic(115),
    to_slogic(118),
    to_slogic(118),
    to_slogic(134),
    to_slogic(152),
    to_slogic(187),
    to_slogic(169),
    to_slogic(165),
    to_slogic(151),
    to_slogic(146),
    to_slogic(146),
    to_slogic(133),
    to_slogic(134),
    to_slogic(128),
    to_slogic(117),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(56),
    to_slogic(56),
    to_slogic(70),
    to_slogic(70),
    to_slogic(64),
    to_slogic(62),
    to_slogic(44),
    to_slogic(56),
    to_slogic(36),
    to_slogic(83),
    to_slogic(162),
    to_slogic(149),
    to_slogic(139),
    to_slogic(109),
    to_slogic(40),
    to_slogic(69),
    to_slogic(118),
    to_slogic(152),
    to_slogic(144),
    to_slogic(143),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(143),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(139),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(132),
    to_slogic(137),
    to_slogic(166),
    to_slogic(183),
    to_slogic(191),
    to_slogic(197),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(204),
    to_slogic(81),
    to_slogic(82),
    to_slogic(75),
    to_slogic(81),
    to_slogic(76),
    to_slogic(76),
    to_slogic(70),
    to_slogic(62),
    to_slogic(70),
    to_slogic(76),
    to_slogic(75),
    to_slogic(92),
    to_slogic(126),
    to_slogic(137),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(165),
    to_slogic(151),
    to_slogic(139),
    to_slogic(121),
    to_slogic(89),
    to_slogic(70),
    to_slogic(81),
    to_slogic(82),
    to_slogic(99),
    to_slogic(92),
    to_slogic(118),
    to_slogic(110),
    to_slogic(119),
    to_slogic(88),
    to_slogic(64),
    to_slogic(50),
    to_slogic(88),
    to_slogic(82),
    to_slogic(75),
    to_slogic(50),
    to_slogic(44),
    to_slogic(107),
    to_slogic(102),
    to_slogic(71),
    to_slogic(84),
    to_slogic(78),
    to_slogic(78),
    to_slogic(58),
    to_slogic(122),
    to_slogic(84),
    to_slogic(117),
    to_slogic(109),
    to_slogic(145),
    to_slogic(107),
    to_slogic(130),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(64),
    to_slogic(152),
    to_slogic(124),
    to_slogic(64),
    to_slogic(33),
    to_slogic(36),
    to_slogic(81),
    to_slogic(95),
    to_slogic(71),
    to_slogic(40),
    to_slogic(83),
    to_slogic(87),
    to_slogic(109),
    to_slogic(110),
    to_slogic(133),
    to_slogic(118),
    to_slogic(107),
    to_slogic(117),
    to_slogic(143),
    to_slogic(196),
    to_slogic(102),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(68),
    to_slogic(68),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(83),
    to_slogic(109),
    to_slogic(89),
    to_slogic(82),
    to_slogic(115),
    to_slogic(115),
    to_slogic(115),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(134),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(151),
    to_slogic(152),
    to_slogic(149),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(149),
    to_slogic(149),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(134),
    to_slogic(126),
    to_slogic(134),
    to_slogic(161),
    to_slogic(179),
    to_slogic(185),
    to_slogic(187),
    to_slogic(172),
    to_slogic(157),
    to_slogic(151),
    to_slogic(146),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(128),
    to_slogic(83),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(82),
    to_slogic(75),
    to_slogic(70),
    to_slogic(62),
    to_slogic(49),
    to_slogic(44),
    to_slogic(36),
    to_slogic(69),
    to_slogic(158),
    to_slogic(149),
    to_slogic(139),
    to_slogic(109),
    to_slogic(56),
    to_slogic(64),
    to_slogic(130),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(150),
    to_slogic(156),
    to_slogic(158),
    to_slogic(155),
    to_slogic(158),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(151),
    to_slogic(150),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(143),
    to_slogic(166),
    to_slogic(191),
    to_slogic(196),
    to_slogic(197),
    to_slogic(196),
    to_slogic(197),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(81),
    to_slogic(75),
    to_slogic(76),
    to_slogic(76),
    to_slogic(75),
    to_slogic(75),
    to_slogic(76),
    to_slogic(70),
    to_slogic(70),
    to_slogic(76),
    to_slogic(82),
    to_slogic(96),
    to_slogic(128),
    to_slogic(146),
    to_slogic(152),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(172),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(82),
    to_slogic(76),
    to_slogic(81),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(102),
    to_slogic(110),
    to_slogic(124),
    to_slogic(110),
    to_slogic(50),
    to_slogic(46),
    to_slogic(84),
    to_slogic(76),
    to_slogic(65),
    to_slogic(50),
    to_slogic(97),
    to_slogic(113),
    to_slogic(56),
    to_slogic(56),
    to_slogic(76),
    to_slogic(76),
    to_slogic(91),
    to_slogic(97),
    to_slogic(109),
    to_slogic(97),
    to_slogic(117),
    to_slogic(91),
    to_slogic(130),
    to_slogic(122),
    to_slogic(138),
    to_slogic(71),
    to_slogic(42),
    to_slogic(49),
    to_slogic(64),
    to_slogic(125),
    to_slogic(144),
    to_slogic(75),
    to_slogic(40),
    to_slogic(49),
    to_slogic(81),
    to_slogic(56),
    to_slogic(68),
    to_slogic(87),
    to_slogic(101),
    to_slogic(110),
    to_slogic(133),
    to_slogic(165),
    to_slogic(149),
    to_slogic(109),
    to_slogic(101),
    to_slogic(120),
    to_slogic(176),
    to_slogic(171),
    to_slogic(56),
    to_slogic(42),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(83),
    to_slogic(109),
    to_slogic(92),
    to_slogic(97),
    to_slogic(99),
    to_slogic(115),
    to_slogic(121),
    to_slogic(118),
    to_slogic(121),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(142),
    to_slogic(144),
    to_slogic(142),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(152),
    to_slogic(149),
    to_slogic(144),
    to_slogic(142),
    to_slogic(134),
    to_slogic(134),
    to_slogic(146),
    to_slogic(162),
    to_slogic(149),
    to_slogic(151),
    to_slogic(187),
    to_slogic(195),
    to_slogic(195),
    to_slogic(187),
    to_slogic(165),
    to_slogic(155),
    to_slogic(149),
    to_slogic(146),
    to_slogic(146),
    to_slogic(134),
    to_slogic(133),
    to_slogic(119),
    to_slogic(64),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(88),
    to_slogic(70),
    to_slogic(82),
    to_slogic(62),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(63),
    to_slogic(144),
    to_slogic(165),
    to_slogic(125),
    to_slogic(101),
    to_slogic(69),
    to_slogic(92),
    to_slogic(137),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(156),
    to_slogic(158),
    to_slogic(155),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(155),
    to_slogic(152),
    to_slogic(149),
    to_slogic(150),
    to_slogic(151),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(150),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(130),
    to_slogic(143),
    to_slogic(178),
    to_slogic(191),
    to_slogic(191),
    to_slogic(196),
    to_slogic(197),
    to_slogic(197),
    to_slogic(205),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(81),
    to_slogic(76),
    to_slogic(76),
    to_slogic(70),
    to_slogic(62),
    to_slogic(62),
    to_slogic(92),
    to_slogic(102),
    to_slogic(128),
    to_slogic(146),
    to_slogic(152),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(152),
    to_slogic(135),
    to_slogic(121),
    to_slogic(89),
    to_slogic(77),
    to_slogic(82),
    to_slogic(82),
    to_slogic(99),
    to_slogic(92),
    to_slogic(109),
    to_slogic(124),
    to_slogic(142),
    to_slogic(128),
    to_slogic(56),
    to_slogic(50),
    to_slogic(84),
    to_slogic(71),
    to_slogic(78),
    to_slogic(91),
    to_slogic(120),
    to_slogic(71),
    to_slogic(50),
    to_slogic(50),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(97),
    to_slogic(107),
    to_slogic(107),
    to_slogic(122),
    to_slogic(84),
    to_slogic(130),
    to_slogic(115),
    to_slogic(138),
    to_slogic(115),
    to_slogic(56),
    to_slogic(64),
    to_slogic(63),
    to_slogic(109),
    to_slogic(101),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(42),
    to_slogic(50),
    to_slogic(109),
    to_slogic(126),
    to_slogic(126),
    to_slogic(155),
    to_slogic(165),
    to_slogic(176),
    to_slogic(102),
    to_slogic(96),
    to_slogic(120),
    to_slogic(165),
    to_slogic(189),
    to_slogic(88),
    to_slogic(42),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(46),
    to_slogic(46),
    to_slogic(83),
    to_slogic(109),
    to_slogic(92),
    to_slogic(89),
    to_slogic(102),
    to_slogic(115),
    to_slogic(118),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(151),
    to_slogic(149),
    to_slogic(152),
    to_slogic(146),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(162),
    to_slogic(187),
    to_slogic(172),
    to_slogic(157),
    to_slogic(187),
    to_slogic(195),
    to_slogic(195),
    to_slogic(187),
    to_slogic(165),
    to_slogic(155),
    to_slogic(149),
    to_slogic(146),
    to_slogic(134),
    to_slogic(133),
    to_slogic(128),
    to_slogic(96),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(68),
    to_slogic(56),
    to_slogic(94),
    to_slogic(64),
    to_slogic(75),
    to_slogic(63),
    to_slogic(62),
    to_slogic(56),
    to_slogic(44),
    to_slogic(46),
    to_slogic(141),
    to_slogic(158),
    to_slogic(132),
    to_slogic(101),
    to_slogic(75),
    to_slogic(110),
    to_slogic(137),
    to_slogic(144),
    to_slogic(152),
    to_slogic(150),
    to_slogic(158),
    to_slogic(155),
    to_slogic(158),
    to_slogic(155),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(143),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(143),
    to_slogic(151),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(130),
    to_slogic(137),
    to_slogic(156),
    to_slogic(184),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(75),
    to_slogic(76),
    to_slogic(70),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(62),
    to_slogic(62),
    to_slogic(62),
    to_slogic(82),
    to_slogic(101),
    to_slogic(133),
    to_slogic(149),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(172),
    to_slogic(152),
    to_slogic(143),
    to_slogic(115),
    to_slogic(92),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(92),
    to_slogic(99),
    to_slogic(103),
    to_slogic(142),
    to_slogic(133),
    to_slogic(96),
    to_slogic(69),
    to_slogic(56),
    to_slogic(82),
    to_slogic(76),
    to_slogic(115),
    to_slogic(113),
    to_slogic(71),
    to_slogic(56),
    to_slogic(44),
    to_slogic(50),
    to_slogic(65),
    to_slogic(71),
    to_slogic(65),
    to_slogic(84),
    to_slogic(78),
    to_slogic(97),
    to_slogic(107),
    to_slogic(91),
    to_slogic(97),
    to_slogic(115),
    to_slogic(130),
    to_slogic(126),
    to_slogic(83),
    to_slogic(75),
    to_slogic(88),
    to_slogic(96),
    to_slogic(87),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(42),
    to_slogic(81),
    to_slogic(152),
    to_slogic(141),
    to_slogic(162),
    to_slogic(165),
    to_slogic(176),
    to_slogic(130),
    to_slogic(96),
    to_slogic(82),
    to_slogic(118),
    to_slogic(189),
    to_slogic(102),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(75),
    to_slogic(109),
    to_slogic(103),
    to_slogic(99),
    to_slogic(115),
    to_slogic(115),
    to_slogic(124),
    to_slogic(130),
    to_slogic(118),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(149),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(149),
    to_slogic(151),
    to_slogic(152),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(172),
    to_slogic(200),
    to_slogic(193),
    to_slogic(169),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(187),
    to_slogic(165),
    to_slogic(151),
    to_slogic(146),
    to_slogic(146),
    to_slogic(142),
    to_slogic(133),
    to_slogic(128),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(69),
    to_slogic(64),
    to_slogic(92),
    to_slogic(64),
    to_slogic(70),
    to_slogic(62),
    to_slogic(62),
    to_slogic(44),
    to_slogic(44),
    to_slogic(46),
    to_slogic(118),
    to_slogic(165),
    to_slogic(139),
    to_slogic(101),
    to_slogic(96),
    to_slogic(118),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(151),
    to_slogic(150),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(150),
    to_slogic(144),
    to_slogic(144),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(130),
    to_slogic(132),
    to_slogic(158),
    to_slogic(183),
    to_slogic(191),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(205),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(204),
    to_slogic(213),
    to_slogic(75),
    to_slogic(70),
    to_slogic(70),
    to_slogic(76),
    to_slogic(70),
    to_slogic(76),
    to_slogic(70),
    to_slogic(62),
    to_slogic(56),
    to_slogic(76),
    to_slogic(82),
    to_slogic(109),
    to_slogic(127),
    to_slogic(146),
    to_slogic(152),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(156),
    to_slogic(135),
    to_slogic(121),
    to_slogic(89),
    to_slogic(62),
    to_slogic(76),
    to_slogic(89),
    to_slogic(99),
    to_slogic(102),
    to_slogic(128),
    to_slogic(133),
    to_slogic(117),
    to_slogic(110),
    to_slogic(63),
    to_slogic(63),
    to_slogic(78),
    to_slogic(118),
    to_slogic(113),
    to_slogic(50),
    to_slogic(63),
    to_slogic(71),
    to_slogic(63),
    to_slogic(56),
    to_slogic(76),
    to_slogic(65),
    to_slogic(71),
    to_slogic(76),
    to_slogic(76),
    to_slogic(84),
    to_slogic(109),
    to_slogic(76),
    to_slogic(91),
    to_slogic(122),
    to_slogic(122),
    to_slogic(127),
    to_slogic(91),
    to_slogic(75),
    to_slogic(121),
    to_slogic(81),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(63),
    to_slogic(75),
    to_slogic(120),
    to_slogic(149),
    to_slogic(157),
    to_slogic(165),
    to_slogic(191),
    to_slogic(171),
    to_slogic(101),
    to_slogic(92),
    to_slogic(91),
    to_slogic(149),
    to_slogic(130),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(62),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(70),
    to_slogic(109),
    to_slogic(101),
    to_slogic(89),
    to_slogic(102),
    to_slogic(115),
    to_slogic(118),
    to_slogic(118),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(118),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(149),
    to_slogic(146),
    to_slogic(146),
    to_slogic(151),
    to_slogic(152),
    to_slogic(146),
    to_slogic(146),
    to_slogic(151),
    to_slogic(146),
    to_slogic(151),
    to_slogic(149),
    to_slogic(162),
    to_slogic(176),
    to_slogic(204),
    to_slogic(195),
    to_slogic(177),
    to_slogic(193),
    to_slogic(200),
    to_slogic(195),
    to_slogic(187),
    to_slogic(165),
    to_slogic(149),
    to_slogic(146),
    to_slogic(149),
    to_slogic(139),
    to_slogic(133),
    to_slogic(101),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(64),
    to_slogic(63),
    to_slogic(64),
    to_slogic(82),
    to_slogic(70),
    to_slogic(75),
    to_slogic(62),
    to_slogic(62),
    to_slogic(49),
    to_slogic(33),
    to_slogic(44),
    to_slogic(109),
    to_slogic(158),
    to_slogic(130),
    to_slogic(101),
    to_slogic(109),
    to_slogic(118),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(150),
    to_slogic(158),
    to_slogic(150),
    to_slogic(156),
    to_slogic(155),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(137),
    to_slogic(130),
    to_slogic(137),
    to_slogic(172),
    to_slogic(183),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(197),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(76),
    to_slogic(70),
    to_slogic(76),
    to_slogic(62),
    to_slogic(76),
    to_slogic(62),
    to_slogic(76),
    to_slogic(63),
    to_slogic(62),
    to_slogic(70),
    to_slogic(82),
    to_slogic(96),
    to_slogic(128),
    to_slogic(146),
    to_slogic(151),
    to_slogic(162),
    to_slogic(157),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(165),
    to_slogic(157),
    to_slogic(143),
    to_slogic(115),
    to_slogic(89),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(82),
    to_slogic(117),
    to_slogic(133),
    to_slogic(110),
    to_slogic(128),
    to_slogic(96),
    to_slogic(63),
    to_slogic(69),
    to_slogic(102),
    to_slogic(120),
    to_slogic(89),
    to_slogic(42),
    to_slogic(56),
    to_slogic(71),
    to_slogic(71),
    to_slogic(58),
    to_slogic(71),
    to_slogic(56),
    to_slogic(83),
    to_slogic(65),
    to_slogic(76),
    to_slogic(71),
    to_slogic(115),
    to_slogic(58),
    to_slogic(78),
    to_slogic(120),
    to_slogic(120),
    to_slogic(115),
    to_slogic(120),
    to_slogic(95),
    to_slogic(130),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(69),
    to_slogic(81),
    to_slogic(101),
    to_slogic(109),
    to_slogic(141),
    to_slogic(162),
    to_slogic(177),
    to_slogic(189),
    to_slogic(118),
    to_slogic(94),
    to_slogic(92),
    to_slogic(132),
    to_slogic(156),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(75),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(64),
    to_slogic(96),
    to_slogic(110),
    to_slogic(92),
    to_slogic(99),
    to_slogic(115),
    to_slogic(115),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(142),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(146),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(162),
    to_slogic(187),
    to_slogic(211),
    to_slogic(200),
    to_slogic(169),
    to_slogic(179),
    to_slogic(204),
    to_slogic(195),
    to_slogic(187),
    to_slogic(165),
    to_slogic(146),
    to_slogic(146),
    to_slogic(134),
    to_slogic(134),
    to_slogic(127),
    to_slogic(75),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(75),
    to_slogic(82),
    to_slogic(70),
    to_slogic(64),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(46),
    to_slogic(109),
    to_slogic(165),
    to_slogic(125),
    to_slogic(110),
    to_slogic(118),
    to_slogic(130),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(149),
    to_slogic(155),
    to_slogic(155),
    to_slogic(150),
    to_slogic(151),
    to_slogic(150),
    to_slogic(149),
    to_slogic(144),
    to_slogic(150),
    to_slogic(149),
    to_slogic(144),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(130),
    to_slogic(132),
    to_slogic(130),
    to_slogic(130),
    to_slogic(166),
    to_slogic(184),
    to_slogic(196),
    to_slogic(196),
    to_slogic(197),
    to_slogic(205),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(204),
    to_slogic(213),
    to_slogic(70),
    to_slogic(70),
    to_slogic(62),
    to_slogic(70),
    to_slogic(63),
    to_slogic(70),
    to_slogic(63),
    to_slogic(62),
    to_slogic(62),
    to_slogic(76),
    to_slogic(75),
    to_slogic(96),
    to_slogic(128),
    to_slogic(139),
    to_slogic(155),
    to_slogic(157),
    to_slogic(173),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(151),
    to_slogic(143),
    to_slogic(121),
    to_slogic(81),
    to_slogic(62),
    to_slogic(81),
    to_slogic(82),
    to_slogic(110),
    to_slogic(142),
    to_slogic(103),
    to_slogic(102),
    to_slogic(127),
    to_slogic(88),
    to_slogic(69),
    to_slogic(82),
    to_slogic(89),
    to_slogic(107),
    to_slogic(71),
    to_slogic(50),
    to_slogic(56),
    to_slogic(71),
    to_slogic(58),
    to_slogic(71),
    to_slogic(71),
    to_slogic(71),
    to_slogic(83),
    to_slogic(71),
    to_slogic(65),
    to_slogic(71),
    to_slogic(89),
    to_slogic(89),
    to_slogic(58),
    to_slogic(76),
    to_slogic(130),
    to_slogic(117),
    to_slogic(130),
    to_slogic(143),
    to_slogic(82),
    to_slogic(33),
    to_slogic(49),
    to_slogic(75),
    to_slogic(120),
    to_slogic(126),
    to_slogic(109),
    to_slogic(117),
    to_slogic(148),
    to_slogic(170),
    to_slogic(191),
    to_slogic(130),
    to_slogic(94),
    to_slogic(92),
    to_slogic(109),
    to_slogic(166),
    to_slogic(64),
    to_slogic(40),
    to_slogic(40),
    to_slogic(75),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(62),
    to_slogic(64),
    to_slogic(64),
    to_slogic(44),
    to_slogic(33),
    to_slogic(63),
    to_slogic(101),
    to_slogic(101),
    to_slogic(82),
    to_slogic(89),
    to_slogic(115),
    to_slogic(115),
    to_slogic(118),
    to_slogic(124),
    to_slogic(121),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(146),
    to_slogic(149),
    to_slogic(151),
    to_slogic(157),
    to_slogic(161),
    to_slogic(187),
    to_slogic(200),
    to_slogic(204),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(193),
    to_slogic(187),
    to_slogic(165),
    to_slogic(142),
    to_slogic(134),
    to_slogic(146),
    to_slogic(134),
    to_slogic(117),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(42),
    to_slogic(56),
    to_slogic(56),
    to_slogic(69),
    to_slogic(75),
    to_slogic(82),
    to_slogic(70),
    to_slogic(70),
    to_slogic(64),
    to_slogic(64),
    to_slogic(49),
    to_slogic(33),
    to_slogic(44),
    to_slogic(91),
    to_slogic(158),
    to_slogic(125),
    to_slogic(109),
    to_slogic(120),
    to_slogic(135),
    to_slogic(144),
    to_slogic(152),
    to_slogic(150),
    to_slogic(158),
    to_slogic(150),
    to_slogic(156),
    to_slogic(158),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(143),
    to_slogic(149),
    to_slogic(144),
    to_slogic(150),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(130),
    to_slogic(130),
    to_slogic(137),
    to_slogic(178),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(205),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(70),
    to_slogic(63),
    to_slogic(62),
    to_slogic(62),
    to_slogic(70),
    to_slogic(70),
    to_slogic(62),
    to_slogic(76),
    to_slogic(62),
    to_slogic(70),
    to_slogic(82),
    to_slogic(96),
    to_slogic(127),
    to_slogic(146),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(157),
    to_slogic(135),
    to_slogic(121),
    to_slogic(82),
    to_slogic(76),
    to_slogic(77),
    to_slogic(87),
    to_slogic(133),
    to_slogic(110),
    to_slogic(102),
    to_slogic(102),
    to_slogic(121),
    to_slogic(81),
    to_slogic(69),
    to_slogic(50),
    to_slogic(89),
    to_slogic(102),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(71),
    to_slogic(58),
    to_slogic(76),
    to_slogic(71),
    to_slogic(91),
    to_slogic(84),
    to_slogic(89),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(84),
    to_slogic(84),
    to_slogic(58),
    to_slogic(89),
    to_slogic(115),
    to_slogic(120),
    to_slogic(138),
    to_slogic(71),
    to_slogic(42),
    to_slogic(56),
    to_slogic(110),
    to_slogic(133),
    to_slogic(171),
    to_slogic(181),
    to_slogic(166),
    to_slogic(191),
    to_slogic(189),
    to_slogic(156),
    to_slogic(94),
    to_slogic(96),
    to_slogic(107),
    to_slogic(153),
    to_slogic(102),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(88),
    to_slogic(62),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(70),
    to_slogic(44),
    to_slogic(44),
    to_slogic(63),
    to_slogic(96),
    to_slogic(96),
    to_slogic(92),
    to_slogic(97),
    to_slogic(99),
    to_slogic(115),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(146),
    to_slogic(157),
    to_slogic(162),
    to_slogic(177),
    to_slogic(173),
    to_slogic(161),
    to_slogic(151),
    to_slogic(162),
    to_slogic(151),
    to_slogic(128),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(75),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(75),
    to_slogic(82),
    to_slogic(64),
    to_slogic(75),
    to_slogic(70),
    to_slogic(62),
    to_slogic(56),
    to_slogic(33),
    to_slogic(36),
    to_slogic(87),
    to_slogic(158),
    to_slogic(141),
    to_slogic(119),
    to_slogic(118),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(149),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(155),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(143),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(139),
    to_slogic(139),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(176),
    to_slogic(183),
    to_slogic(196),
    to_slogic(203),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(63),
    to_slogic(62),
    to_slogic(62),
    to_slogic(62),
    to_slogic(62),
    to_slogic(70),
    to_slogic(63),
    to_slogic(62),
    to_slogic(56),
    to_slogic(70),
    to_slogic(81),
    to_slogic(96),
    to_slogic(128),
    to_slogic(146),
    to_slogic(155),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(151),
    to_slogic(135),
    to_slogic(121),
    to_slogic(81),
    to_slogic(70),
    to_slogic(77),
    to_slogic(117),
    to_slogic(121),
    to_slogic(92),
    to_slogic(99),
    to_slogic(110),
    to_slogic(142),
    to_slogic(81),
    to_slogic(50),
    to_slogic(46),
    to_slogic(89),
    to_slogic(102),
    to_slogic(65),
    to_slogic(63),
    to_slogic(63),
    to_slogic(65),
    to_slogic(56),
    to_slogic(58),
    to_slogic(65),
    to_slogic(91),
    to_slogic(107),
    to_slogic(91),
    to_slogic(97),
    to_slogic(89),
    to_slogic(76),
    to_slogic(71),
    to_slogic(97),
    to_slogic(84),
    to_slogic(58),
    to_slogic(91),
    to_slogic(109),
    to_slogic(122),
    to_slogic(115),
    to_slogic(76),
    to_slogic(102),
    to_slogic(121),
    to_slogic(113),
    to_slogic(170),
    to_slogic(197),
    to_slogic(204),
    to_slogic(204),
    to_slogic(166),
    to_slogic(102),
    to_slogic(94),
    to_slogic(96),
    to_slogic(143),
    to_slogic(143),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(75),
    to_slogic(62),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(75),
    to_slogic(70),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(91),
    to_slogic(96),
    to_slogic(82),
    to_slogic(81),
    to_slogic(99),
    to_slogic(115),
    to_slogic(115),
    to_slogic(121),
    to_slogic(130),
    to_slogic(124),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(121),
    to_slogic(115),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(134),
    to_slogic(135),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(134),
    to_slogic(118),
    to_slogic(121),
    to_slogic(118),
    to_slogic(134),
    to_slogic(134),
    to_slogic(146),
    to_slogic(134),
    to_slogic(118),
    to_slogic(126),
    to_slogic(134),
    to_slogic(102),
    to_slogic(118),
    to_slogic(134),
    to_slogic(146),
    to_slogic(119),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(63),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(33),
    to_slogic(44),
    to_slogic(75),
    to_slogic(149),
    to_slogic(133),
    to_slogic(120),
    to_slogic(130),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(150),
    to_slogic(158),
    to_slogic(149),
    to_slogic(158),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(144),
    to_slogic(144),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(130),
    to_slogic(125),
    to_slogic(143),
    to_slogic(172),
    to_slogic(191),
    to_slogic(197),
    to_slogic(205),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(62),
    to_slogic(70),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(76),
    to_slogic(82),
    to_slogic(102),
    to_slogic(127),
    to_slogic(146),
    to_slogic(151),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(172),
    to_slogic(157),
    to_slogic(135),
    to_slogic(121),
    to_slogic(82),
    to_slogic(77),
    to_slogic(110),
    to_slogic(133),
    to_slogic(92),
    to_slogic(82),
    to_slogic(110),
    to_slogic(133),
    to_slogic(141),
    to_slogic(69),
    to_slogic(50),
    to_slogic(69),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(65),
    to_slogic(63),
    to_slogic(83),
    to_slogic(65),
    to_slogic(44),
    to_slogic(58),
    to_slogic(97),
    to_slogic(130),
    to_slogic(107),
    to_slogic(97),
    to_slogic(97),
    to_slogic(84),
    to_slogic(76),
    to_slogic(71),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(71),
    to_slogic(107),
    to_slogic(76),
    to_slogic(107),
    to_slogic(148),
    to_slogic(134),
    to_slogic(143),
    to_slogic(193),
    to_slogic(197),
    to_slogic(204),
    to_slogic(189),
    to_slogic(101),
    to_slogic(109),
    to_slogic(96),
    to_slogic(119),
    to_slogic(171),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(62),
    to_slogic(70),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(75),
    to_slogic(49),
    to_slogic(36),
    to_slogic(56),
    to_slogic(91),
    to_slogic(82),
    to_slogic(92),
    to_slogic(76),
    to_slogic(97),
    to_slogic(115),
    to_slogic(115),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(121),
    to_slogic(124),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(135),
    to_slogic(97),
    to_slogic(81),
    to_slogic(81),
    to_slogic(97),
    to_slogic(97),
    to_slogic(109),
    to_slogic(115),
    to_slogic(97),
    to_slogic(115),
    to_slogic(99),
    to_slogic(97),
    to_slogic(97),
    to_slogic(97),
    to_slogic(97),
    to_slogic(99),
    to_slogic(118),
    to_slogic(121),
    to_slogic(121),
    to_slogic(97),
    to_slogic(76),
    to_slogic(99),
    to_slogic(109),
    to_slogic(118),
    to_slogic(128),
    to_slogic(146),
    to_slogic(139),
    to_slogic(82),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(63),
    to_slogic(75),
    to_slogic(70),
    to_slogic(75),
    to_slogic(75),
    to_slogic(56),
    to_slogic(62),
    to_slogic(70),
    to_slogic(44),
    to_slogic(36),
    to_slogic(64),
    to_slogic(143),
    to_slogic(141),
    to_slogic(137),
    to_slogic(137),
    to_slogic(144),
    to_slogic(151),
    to_slogic(143),
    to_slogic(149),
    to_slogic(158),
    to_slogic(158),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(130),
    to_slogic(132),
    to_slogic(130),
    to_slogic(143),
    to_slogic(176),
    to_slogic(191),
    to_slogic(203),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(63),
    to_slogic(63),
    to_slogic(62),
    to_slogic(63),
    to_slogic(62),
    to_slogic(82),
    to_slogic(82),
    to_slogic(101),
    to_slogic(128),
    to_slogic(151),
    to_slogic(157),
    to_slogic(162),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(165),
    to_slogic(152),
    to_slogic(135),
    to_slogic(116),
    to_slogic(82),
    to_slogic(96),
    to_slogic(142),
    to_slogic(102),
    to_slogic(82),
    to_slogic(99),
    to_slogic(128),
    to_slogic(142),
    to_slogic(121),
    to_slogic(69),
    to_slogic(65),
    to_slogic(71),
    to_slogic(56),
    to_slogic(42),
    to_slogic(56),
    to_slogic(71),
    to_slogic(68),
    to_slogic(76),
    to_slogic(56),
    to_slogic(76),
    to_slogic(58),
    to_slogic(102),
    to_slogic(130),
    to_slogic(109),
    to_slogic(97),
    to_slogic(103),
    to_slogic(103),
    to_slogic(103),
    to_slogic(84),
    to_slogic(84),
    to_slogic(120),
    to_slogic(115),
    to_slogic(65),
    to_slogic(76),
    to_slogic(65),
    to_slogic(102),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(197),
    to_slogic(214),
    to_slogic(205),
    to_slogic(149),
    to_slogic(94),
    to_slogic(92),
    to_slogic(109),
    to_slogic(170),
    to_slogic(114),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(75),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(83),
    to_slogic(82),
    to_slogic(83),
    to_slogic(81),
    to_slogic(89),
    to_slogic(99),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(134),
    to_slogic(118),
    to_slogic(118),
    to_slogic(115),
    to_slogic(99),
    to_slogic(99),
    to_slogic(97),
    to_slogic(97),
    to_slogic(118),
    to_slogic(118),
    to_slogic(115),
    to_slogic(115),
    to_slogic(115),
    to_slogic(99),
    to_slogic(118),
    to_slogic(118),
    to_slogic(118),
    to_slogic(142),
    to_slogic(124),
    to_slogic(142),
    to_slogic(124),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(144),
    to_slogic(109),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(56),
    to_slogic(56),
    to_slogic(82),
    to_slogic(44),
    to_slogic(46),
    to_slogic(56),
    to_slogic(134),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(143),
    to_slogic(151),
    to_slogic(152),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(158),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(132),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(157),
    to_slogic(183),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(62),
    to_slogic(62),
    to_slogic(62),
    to_slogic(70),
    to_slogic(82),
    to_slogic(87),
    to_slogic(110),
    to_slogic(133),
    to_slogic(146),
    to_slogic(151),
    to_slogic(162),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(178),
    to_slogic(165),
    to_slogic(151),
    to_slogic(139),
    to_slogic(118),
    to_slogic(110),
    to_slogic(152),
    to_slogic(103),
    to_slogic(81),
    to_slogic(82),
    to_slogic(103),
    to_slogic(142),
    to_slogic(128),
    to_slogic(110),
    to_slogic(75),
    to_slogic(69),
    to_slogic(63),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(56),
    to_slogic(76),
    to_slogic(58),
    to_slogic(78),
    to_slogic(58),
    to_slogic(115),
    to_slogic(153),
    to_slogic(97),
    to_slogic(84),
    to_slogic(91),
    to_slogic(97),
    to_slogic(102),
    to_slogic(97),
    to_slogic(89),
    to_slogic(83),
    to_slogic(89),
    to_slogic(91),
    to_slogic(84),
    to_slogic(97),
    to_slogic(133),
    to_slogic(151),
    to_slogic(130),
    to_slogic(126),
    to_slogic(172),
    to_slogic(220),
    to_slogic(176),
    to_slogic(109),
    to_slogic(101),
    to_slogic(107),
    to_slogic(166),
    to_slogic(156),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(75),
    to_slogic(64),
    to_slogic(44),
    to_slogic(56),
    to_slogic(83),
    to_slogic(75),
    to_slogic(83),
    to_slogic(75),
    to_slogic(89),
    to_slogic(100),
    to_slogic(115),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(118),
    to_slogic(121),
    to_slogic(130),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(139),
    to_slogic(144),
    to_slogic(134),
    to_slogic(130),
    to_slogic(124),
    to_slogic(121),
    to_slogic(118),
    to_slogic(118),
    to_slogic(118),
    to_slogic(118),
    to_slogic(134),
    to_slogic(126),
    to_slogic(142),
    to_slogic(151),
    to_slogic(154),
    to_slogic(161),
    to_slogic(161),
    to_slogic(175),
    to_slogic(183),
    to_slogic(179),
    to_slogic(161),
    to_slogic(127),
    to_slogic(142),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(133),
    to_slogic(75),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(63),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(56),
    to_slogic(62),
    to_slogic(82),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(125),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(143),
    to_slogic(150),
    to_slogic(158),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(139),
    to_slogic(130),
    to_slogic(125),
    to_slogic(150),
    to_slogic(183),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(62),
    to_slogic(62),
    to_slogic(56),
    to_slogic(63),
    to_slogic(82),
    to_slogic(92),
    to_slogic(101),
    to_slogic(128),
    to_slogic(139),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(173),
    to_slogic(165),
    to_slogic(157),
    to_slogic(142),
    to_slogic(124),
    to_slogic(141),
    to_slogic(101),
    to_slogic(76),
    to_slogic(77),
    to_slogic(81),
    to_slogic(133),
    to_slogic(133),
    to_slogic(110),
    to_slogic(103),
    to_slogic(81),
    to_slogic(65),
    to_slogic(81),
    to_slogic(84),
    to_slogic(56),
    to_slogic(40),
    to_slogic(44),
    to_slogic(56),
    to_slogic(89),
    to_slogic(56),
    to_slogic(84),
    to_slogic(58),
    to_slogic(117),
    to_slogic(153),
    to_slogic(97),
    to_slogic(58),
    to_slogic(91),
    to_slogic(107),
    to_slogic(109),
    to_slogic(91),
    to_slogic(91),
    to_slogic(71),
    to_slogic(65),
    to_slogic(97),
    to_slogic(107),
    to_slogic(130),
    to_slogic(133),
    to_slogic(146),
    to_slogic(130),
    to_slogic(126),
    to_slogic(157),
    to_slogic(196),
    to_slogic(118),
    to_slogic(101),
    to_slogic(128),
    to_slogic(166),
    to_slogic(171),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(70),
    to_slogic(44),
    to_slogic(62),
    to_slogic(82),
    to_slogic(70),
    to_slogic(82),
    to_slogic(70),
    to_slogic(81),
    to_slogic(99),
    to_slogic(109),
    to_slogic(115),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(124),
    to_slogic(118),
    to_slogic(134),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(142),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(139),
    to_slogic(134),
    to_slogic(130),
    to_slogic(118),
    to_slogic(121),
    to_slogic(124),
    to_slogic(118),
    to_slogic(118),
    to_slogic(118),
    to_slogic(134),
    to_slogic(142),
    to_slogic(157),
    to_slogic(172),
    to_slogic(169),
    to_slogic(169),
    to_slogic(177),
    to_slogic(183),
    to_slogic(187),
    to_slogic(154),
    to_slogic(142),
    to_slogic(134),
    to_slogic(152),
    to_slogic(146),
    to_slogic(137),
    to_slogic(96),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(62),
    to_slogic(83),
    to_slogic(75),
    to_slogic(75),
    to_slogic(76),
    to_slogic(49),
    to_slogic(70),
    to_slogic(82),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(120),
    to_slogic(165),
    to_slogic(139),
    to_slogic(152),
    to_slogic(150),
    to_slogic(151),
    to_slogic(150),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(158),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(132),
    to_slogic(130),
    to_slogic(132),
    to_slogic(124),
    to_slogic(158),
    to_slogic(183),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(83),
    to_slogic(92),
    to_slogic(96),
    to_slogic(127),
    to_slogic(146),
    to_slogic(157),
    to_slogic(151),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(173),
    to_slogic(169),
    to_slogic(155),
    to_slogic(142),
    to_slogic(102),
    to_slogic(63),
    to_slogic(76),
    to_slogic(82),
    to_slogic(110),
    to_slogic(142),
    to_slogic(110),
    to_slogic(110),
    to_slogic(96),
    to_slogic(69),
    to_slogic(71),
    to_slogic(115),
    to_slogic(89),
    to_slogic(49),
    to_slogic(42),
    to_slogic(42),
    to_slogic(83),
    to_slogic(78),
    to_slogic(76),
    to_slogic(76),
    to_slogic(78),
    to_slogic(130),
    to_slogic(145),
    to_slogic(117),
    to_slogic(58),
    to_slogic(78),
    to_slogic(84),
    to_slogic(91),
    to_slogic(115),
    to_slogic(107),
    to_slogic(84),
    to_slogic(78),
    to_slogic(89),
    to_slogic(103),
    to_slogic(132),
    to_slogic(141),
    to_slogic(152),
    to_slogic(124),
    to_slogic(134),
    to_slogic(196),
    to_slogic(149),
    to_slogic(101),
    to_slogic(130),
    to_slogic(166),
    to_slogic(158),
    to_slogic(88),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(63),
    to_slogic(64),
    to_slogic(70),
    to_slogic(49),
    to_slogic(49),
    to_slogic(75),
    to_slogic(64),
    to_slogic(82),
    to_slogic(70),
    to_slogic(75),
    to_slogic(97),
    to_slogic(99),
    to_slogic(109),
    to_slogic(115),
    to_slogic(115),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(118),
    to_slogic(130),
    to_slogic(124),
    to_slogic(118),
    to_slogic(142),
    to_slogic(142),
    to_slogic(142),
    to_slogic(149),
    to_slogic(151),
    to_slogic(142),
    to_slogic(142),
    to_slogic(151),
    to_slogic(142),
    to_slogic(134),
    to_slogic(146),
    to_slogic(151),
    to_slogic(137),
    to_slogic(128),
    to_slogic(62),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(44),
    to_slogic(70),
    to_slogic(83),
    to_slogic(76),
    to_slogic(82),
    to_slogic(75),
    to_slogic(62),
    to_slogic(64),
    to_slogic(82),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(109),
    to_slogic(162),
    to_slogic(143),
    to_slogic(157),
    to_slogic(157),
    to_slogic(144),
    to_slogic(150),
    to_slogic(156),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(130),
    to_slogic(125),
    to_slogic(125),
    to_slogic(158),
    to_slogic(191),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(82),
    to_slogic(94),
    to_slogic(96),
    to_slogic(126),
    to_slogic(144),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(183),
    to_slogic(172),
    to_slogic(165),
    to_slogic(157),
    to_slogic(146),
    to_slogic(124),
    to_slogic(81),
    to_slogic(63),
    to_slogic(77),
    to_slogic(87),
    to_slogic(142),
    to_slogic(128),
    to_slogic(102),
    to_slogic(110),
    to_slogic(87),
    to_slogic(56),
    to_slogic(65),
    to_slogic(138),
    to_slogic(63),
    to_slogic(42),
    to_slogic(49),
    to_slogic(50),
    to_slogic(97),
    to_slogic(65),
    to_slogic(78),
    to_slogic(84),
    to_slogic(84),
    to_slogic(155),
    to_slogic(122),
    to_slogic(120),
    to_slogic(86),
    to_slogic(78),
    to_slogic(102),
    to_slogic(65),
    to_slogic(97),
    to_slogic(115),
    to_slogic(115),
    to_slogic(109),
    to_slogic(122),
    to_slogic(103),
    to_slogic(143),
    to_slogic(160),
    to_slogic(141),
    to_slogic(126),
    to_slogic(149),
    to_slogic(191),
    to_slogic(120),
    to_slogic(133),
    to_slogic(172),
    to_slogic(191),
    to_slogic(114),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(82),
    to_slogic(75),
    to_slogic(82),
    to_slogic(62),
    to_slogic(70),
    to_slogic(89),
    to_slogic(97),
    to_slogic(109),
    to_slogic(115),
    to_slogic(115),
    to_slogic(115),
    to_slogic(115),
    to_slogic(124),
    to_slogic(121),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(146),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(121),
    to_slogic(126),
    to_slogic(118),
    to_slogic(134),
    to_slogic(142),
    to_slogic(142),
    to_slogic(142),
    to_slogic(142),
    to_slogic(134),
    to_slogic(134),
    to_slogic(142),
    to_slogic(149),
    to_slogic(146),
    to_slogic(146),
    to_slogic(133),
    to_slogic(101),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(70),
    to_slogic(83),
    to_slogic(70),
    to_slogic(82),
    to_slogic(75),
    to_slogic(70),
    to_slogic(62),
    to_slogic(82),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(120),
    to_slogic(158),
    to_slogic(155),
    to_slogic(152),
    to_slogic(150),
    to_slogic(152),
    to_slogic(150),
    to_slogic(150),
    to_slogic(156),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(130),
    to_slogic(119),
    to_slogic(124),
    to_slogic(158),
    to_slogic(197),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(92),
    to_slogic(83),
    to_slogic(92),
    to_slogic(119),
    to_slogic(144),
    to_slogic(152),
    to_slogic(155),
    to_slogic(165),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(173),
    to_slogic(157),
    to_slogic(139),
    to_slogic(109),
    to_slogic(76),
    to_slogic(77),
    to_slogic(64),
    to_slogic(117),
    to_slogic(142),
    to_slogic(103),
    to_slogic(96),
    to_slogic(117),
    to_slogic(69),
    to_slogic(58),
    to_slogic(81),
    to_slogic(143),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(50),
    to_slogic(102),
    to_slogic(65),
    to_slogic(56),
    to_slogic(84),
    to_slogic(91),
    to_slogic(168),
    to_slogic(117),
    to_slogic(78),
    to_slogic(130),
    to_slogic(107),
    to_slogic(122),
    to_slogic(78),
    to_slogic(65),
    to_slogic(84),
    to_slogic(130),
    to_slogic(132),
    to_slogic(113),
    to_slogic(126),
    to_slogic(107),
    to_slogic(155),
    to_slogic(133),
    to_slogic(128),
    to_slogic(143),
    to_slogic(197),
    to_slogic(150),
    to_slogic(162),
    to_slogic(191),
    to_slogic(124),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(64),
    to_slogic(75),
    to_slogic(56),
    to_slogic(49),
    to_slogic(75),
    to_slogic(70),
    to_slogic(82),
    to_slogic(64),
    to_slogic(70),
    to_slogic(76),
    to_slogic(89),
    to_slogic(109),
    to_slogic(97),
    to_slogic(109),
    to_slogic(115),
    to_slogic(121),
    to_slogic(118),
    to_slogic(124),
    to_slogic(124),
    to_slogic(130),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(124),
    to_slogic(134),
    to_slogic(121),
    to_slogic(124),
    to_slogic(115),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(126),
    to_slogic(115),
    to_slogic(118),
    to_slogic(124),
    to_slogic(142),
    to_slogic(151),
    to_slogic(146),
    to_slogic(146),
    to_slogic(144),
    to_slogic(94),
    to_slogic(75),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(44),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(70),
    to_slogic(56),
    to_slogic(82),
    to_slogic(62),
    to_slogic(44),
    to_slogic(56),
    to_slogic(109),
    to_slogic(158),
    to_slogic(152),
    to_slogic(157),
    to_slogic(150),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(158),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(130),
    to_slogic(124),
    to_slogic(125),
    to_slogic(158),
    to_slogic(197),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(223),
    to_slogic(213),
    to_slogic(223),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(70),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(117),
    to_slogic(137),
    to_slogic(144),
    to_slogic(155),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(173),
    to_slogic(165),
    to_slogic(152),
    to_slogic(139),
    to_slogic(121),
    to_slogic(76),
    to_slogic(63),
    to_slogic(77),
    to_slogic(121),
    to_slogic(121),
    to_slogic(103),
    to_slogic(110),
    to_slogic(87),
    to_slogic(50),
    to_slogic(56),
    to_slogic(89),
    to_slogic(127),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(71),
    to_slogic(84),
    to_slogic(56),
    to_slogic(44),
    to_slogic(71),
    to_slogic(109),
    to_slogic(168),
    to_slogic(132),
    to_slogic(76),
    to_slogic(122),
    to_slogic(122),
    to_slogic(122),
    to_slogic(91),
    to_slogic(78),
    to_slogic(78),
    to_slogic(130),
    to_slogic(130),
    to_slogic(115),
    to_slogic(113),
    to_slogic(83),
    to_slogic(127),
    to_slogic(113),
    to_slogic(121),
    to_slogic(162),
    to_slogic(185),
    to_slogic(157),
    to_slogic(177),
    to_slogic(158),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(64),
    to_slogic(82),
    to_slogic(64),
    to_slogic(64),
    to_slogic(70),
    to_slogic(81),
    to_slogic(97),
    to_slogic(97),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(115),
    to_slogic(124),
    to_slogic(124),
    to_slogic(130),
    to_slogic(134),
    to_slogic(134),
    to_slogic(142),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(124),
    to_slogic(118),
    to_slogic(126),
    to_slogic(126),
    to_slogic(134),
    to_slogic(139),
    to_slogic(149),
    to_slogic(151),
    to_slogic(149),
    to_slogic(142),
    to_slogic(137),
    to_slogic(128),
    to_slogic(62),
    to_slogic(64),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(75),
    to_slogic(96),
    to_slogic(76),
    to_slogic(82),
    to_slogic(75),
    to_slogic(70),
    to_slogic(64),
    to_slogic(82),
    to_slogic(62),
    to_slogic(56),
    to_slogic(50),
    to_slogic(109),
    to_slogic(172),
    to_slogic(143),
    to_slogic(157),
    to_slogic(152),
    to_slogic(143),
    to_slogic(158),
    to_slogic(156),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(130),
    to_slogic(130),
    to_slogic(119),
    to_slogic(118),
    to_slogic(158),
    to_slogic(198),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(56),
    to_slogic(44),
    to_slogic(49),
    to_slogic(83),
    to_slogic(94),
    to_slogic(109),
    to_slogic(96),
    to_slogic(126),
    to_slogic(133),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(173),
    to_slogic(157),
    to_slogic(135),
    to_slogic(121),
    to_slogic(82),
    to_slogic(63),
    to_slogic(77),
    to_slogic(121),
    to_slogic(121),
    to_slogic(96),
    to_slogic(96),
    to_slogic(81),
    to_slogic(65),
    to_slogic(56),
    to_slogic(89),
    to_slogic(89),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(71),
    to_slogic(71),
    to_slogic(63),
    to_slogic(58),
    to_slogic(44),
    to_slogic(130),
    to_slogic(155),
    to_slogic(130),
    to_slogic(117),
    to_slogic(97),
    to_slogic(140),
    to_slogic(130),
    to_slogic(107),
    to_slogic(107),
    to_slogic(115),
    to_slogic(91),
    to_slogic(117),
    to_slogic(120),
    to_slogic(88),
    to_slogic(84),
    to_slogic(130),
    to_slogic(107),
    to_slogic(122),
    to_slogic(166),
    to_slogic(191),
    to_slogic(183),
    to_slogic(183),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(64),
    to_slogic(62),
    to_slogic(75),
    to_slogic(81),
    to_slogic(89),
    to_slogic(89),
    to_slogic(97),
    to_slogic(109),
    to_slogic(99),
    to_slogic(115),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(128),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(149),
    to_slogic(149),
    to_slogic(146),
    to_slogic(149),
    to_slogic(149),
    to_slogic(151),
    to_slogic(151),
    to_slogic(146),
    to_slogic(146),
    to_slogic(137),
    to_slogic(92),
    to_slogic(49),
    to_slogic(64),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(75),
    to_slogic(83),
    to_slogic(75),
    to_slogic(94),
    to_slogic(75),
    to_slogic(64),
    to_slogic(62),
    to_slogic(75),
    to_slogic(70),
    to_slogic(49),
    to_slogic(50),
    to_slogic(101),
    to_slogic(167),
    to_slogic(155),
    to_slogic(157),
    to_slogic(143),
    to_slogic(150),
    to_slogic(158),
    to_slogic(150),
    to_slogic(156),
    to_slogic(158),
    to_slogic(156),
    to_slogic(149),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(132),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(124),
    to_slogic(119),
    to_slogic(124),
    to_slogic(158),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(223),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(62),
    to_slogic(92),
    to_slogic(109),
    to_slogic(96),
    to_slogic(109),
    to_slogic(124),
    to_slogic(133),
    to_slogic(144),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(157),
    to_slogic(143),
    to_slogic(115),
    to_slogic(81),
    to_slogic(76),
    to_slogic(64),
    to_slogic(110),
    to_slogic(121),
    to_slogic(103),
    to_slogic(96),
    to_slogic(81),
    to_slogic(63),
    to_slogic(88),
    to_slogic(81),
    to_slogic(68),
    to_slogic(56),
    to_slogic(42),
    to_slogic(42),
    to_slogic(81),
    to_slogic(71),
    to_slogic(56),
    to_slogic(58),
    to_slogic(58),
    to_slogic(113),
    to_slogic(153),
    to_slogic(117),
    to_slogic(115),
    to_slogic(107),
    to_slogic(140),
    to_slogic(138),
    to_slogic(107),
    to_slogic(115),
    to_slogic(91),
    to_slogic(84),
    to_slogic(107),
    to_slogic(127),
    to_slogic(103),
    to_slogic(81),
    to_slogic(120),
    to_slogic(102),
    to_slogic(121),
    to_slogic(185),
    to_slogic(211),
    to_slogic(191),
    to_slogic(88),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(62),
    to_slogic(75),
    to_slogic(56),
    to_slogic(62),
    to_slogic(62),
    to_slogic(76),
    to_slogic(97),
    to_slogic(97),
    to_slogic(97),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(127),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(151),
    to_slogic(161),
    to_slogic(165),
    to_slogic(165),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(151),
    to_slogic(149),
    to_slogic(149),
    to_slogic(146),
    to_slogic(133),
    to_slogic(49),
    to_slogic(62),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(82),
    to_slogic(96),
    to_slogic(70),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(70),
    to_slogic(82),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(101),
    to_slogic(167),
    to_slogic(156),
    to_slogic(165),
    to_slogic(144),
    to_slogic(143),
    to_slogic(158),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(150),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(149),
    to_slogic(143),
    to_slogic(133),
    to_slogic(132),
    to_slogic(132),
    to_slogic(119),
    to_slogic(119),
    to_slogic(120),
    to_slogic(158),
    to_slogic(207),
    to_slogic(213),
    to_slogic(223),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(96),
    to_slogic(102),
    to_slogic(96),
    to_slogic(102),
    to_slogic(118),
    to_slogic(139),
    to_slogic(144),
    to_slogic(152),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(157),
    to_slogic(135),
    to_slogic(121),
    to_slogic(82),
    to_slogic(63),
    to_slogic(77),
    to_slogic(87),
    to_slogic(113),
    to_slogic(110),
    to_slogic(88),
    to_slogic(75),
    to_slogic(75),
    to_slogic(95),
    to_slogic(89),
    to_slogic(63),
    to_slogic(49),
    to_slogic(42),
    to_slogic(42),
    to_slogic(89),
    to_slogic(71),
    to_slogic(44),
    to_slogic(56),
    to_slogic(58),
    to_slogic(97),
    to_slogic(130),
    to_slogic(102),
    to_slogic(109),
    to_slogic(117),
    to_slogic(109),
    to_slogic(140),
    to_slogic(109),
    to_slogic(117),
    to_slogic(97),
    to_slogic(84),
    to_slogic(78),
    to_slogic(127),
    to_slogic(110),
    to_slogic(110),
    to_slogic(122),
    to_slogic(81),
    to_slogic(113),
    to_slogic(144),
    to_slogic(193),
    to_slogic(102),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(62),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(62),
    to_slogic(64),
    to_slogic(49),
    to_slogic(62),
    to_slogic(70),
    to_slogic(56),
    to_slogic(62),
    to_slogic(89),
    to_slogic(97),
    to_slogic(97),
    to_slogic(109),
    to_slogic(115),
    to_slogic(121),
    to_slogic(124),
    to_slogic(134),
    to_slogic(128),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(142),
    to_slogic(146),
    to_slogic(144),
    to_slogic(149),
    to_slogic(149),
    to_slogic(152),
    to_slogic(149),
    to_slogic(151),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(151),
    to_slogic(157),
    to_slogic(151),
    to_slogic(151),
    to_slogic(146),
    to_slogic(152),
    to_slogic(96),
    to_slogic(40),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(82),
    to_slogic(96),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(70),
    to_slogic(75),
    to_slogic(82),
    to_slogic(70),
    to_slogic(63),
    to_slogic(50),
    to_slogic(101),
    to_slogic(172),
    to_slogic(162),
    to_slogic(162),
    to_slogic(143),
    to_slogic(156),
    to_slogic(158),
    to_slogic(156),
    to_slogic(158),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(156),
    to_slogic(149),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(143),
    to_slogic(133),
    to_slogic(149),
    to_slogic(143),
    to_slogic(130),
    to_slogic(130),
    to_slogic(119),
    to_slogic(124),
    to_slogic(166),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(223),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(44),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(46),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(94),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(126),
    to_slogic(133),
    to_slogic(144),
    to_slogic(151),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(172),
    to_slogic(152),
    to_slogic(143),
    to_slogic(115),
    to_slogic(81),
    to_slogic(76),
    to_slogic(70),
    to_slogic(92),
    to_slogic(110),
    to_slogic(96),
    to_slogic(96),
    to_slogic(63),
    to_slogic(75),
    to_slogic(75),
    to_slogic(95),
    to_slogic(63),
    to_slogic(56),
    to_slogic(44),
    to_slogic(42),
    to_slogic(83),
    to_slogic(65),
    to_slogic(49),
    to_slogic(56),
    to_slogic(76),
    to_slogic(97),
    to_slogic(120),
    to_slogic(97),
    to_slogic(78),
    to_slogic(97),
    to_slogic(122),
    to_slogic(122),
    to_slogic(132),
    to_slogic(122),
    to_slogic(117),
    to_slogic(103),
    to_slogic(78),
    to_slogic(130),
    to_slogic(113),
    to_slogic(124),
    to_slogic(126),
    to_slogic(65),
    to_slogic(102),
    to_slogic(133),
    to_slogic(177),
    to_slogic(63),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(75),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(76),
    to_slogic(97),
    to_slogic(97),
    to_slogic(97),
    to_slogic(115),
    to_slogic(121),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(133),
    to_slogic(142),
    to_slogic(146),
    to_slogic(134),
    to_slogic(146),
    to_slogic(149),
    to_slogic(157),
    to_slogic(162),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(157),
    to_slogic(149),
    to_slogic(151),
    to_slogic(139),
    to_slogic(70),
    to_slogic(49),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(64),
    to_slogic(49),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(91),
    to_slogic(96),
    to_slogic(82),
    to_slogic(91),
    to_slogic(82),
    to_slogic(70),
    to_slogic(75),
    to_slogic(75),
    to_slogic(70),
    to_slogic(63),
    to_slogic(49),
    to_slogic(101),
    to_slogic(165),
    to_slogic(156),
    to_slogic(162),
    to_slogic(137),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(156),
    to_slogic(150),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(119),
    to_slogic(119),
    to_slogic(130),
    to_slogic(171),
    to_slogic(213),
    to_slogic(213),
    to_slogic(223),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(198),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(70),
    to_slogic(89),
    to_slogic(96),
    to_slogic(94),
    to_slogic(109),
    to_slogic(126),
    to_slogic(135),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(176),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(165),
    to_slogic(157),
    to_slogic(135),
    to_slogic(121),
    to_slogic(82),
    to_slogic(63),
    to_slogic(77),
    to_slogic(92),
    to_slogic(96),
    to_slogic(96),
    to_slogic(68),
    to_slogic(63),
    to_slogic(56),
    to_slogic(71),
    to_slogic(107),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(50),
    to_slogic(81),
    to_slogic(65),
    to_slogic(50),
    to_slogic(58),
    to_slogic(65),
    to_slogic(102),
    to_slogic(115),
    to_slogic(97),
    to_slogic(56),
    to_slogic(58),
    to_slogic(76),
    to_slogic(122),
    to_slogic(140),
    to_slogic(132),
    to_slogic(122),
    to_slogic(122),
    to_slogic(107),
    to_slogic(122),
    to_slogic(127),
    to_slogic(128),
    to_slogic(141),
    to_slogic(89),
    to_slogic(91),
    to_slogic(91),
    to_slogic(114),
    to_slogic(68),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(56),
    to_slogic(75),
    to_slogic(62),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(76),
    to_slogic(89),
    to_slogic(97),
    to_slogic(99),
    to_slogic(115),
    to_slogic(124),
    to_slogic(126),
    to_slogic(128),
    to_slogic(139),
    to_slogic(134),
    to_slogic(133),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(151),
    to_slogic(151),
    to_slogic(165),
    to_slogic(169),
    to_slogic(162),
    to_slogic(161),
    to_slogic(162),
    to_slogic(165),
    to_slogic(161),
    to_slogic(165),
    to_slogic(169),
    to_slogic(169),
    to_slogic(155),
    to_slogic(149),
    to_slogic(152),
    to_slogic(117),
    to_slogic(49),
    to_slogic(40),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(44),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(96),
    to_slogic(96),
    to_slogic(82),
    to_slogic(91),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(62),
    to_slogic(75),
    to_slogic(49),
    to_slogic(96),
    to_slogic(172),
    to_slogic(162),
    to_slogic(162),
    to_slogic(143),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(158),
    to_slogic(156),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(114),
    to_slogic(119),
    to_slogic(183),
    to_slogic(213),
    to_slogic(223),
    to_slogic(223),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(205),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(205),
    to_slogic(191),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(82),
    to_slogic(92),
    to_slogic(94),
    to_slogic(109),
    to_slogic(126),
    to_slogic(139),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(157),
    to_slogic(135),
    to_slogic(121),
    to_slogic(81),
    to_slogic(63),
    to_slogic(76),
    to_slogic(83),
    to_slogic(110),
    to_slogic(83),
    to_slogic(50),
    to_slogic(56),
    to_slogic(56),
    to_slogic(81),
    to_slogic(107),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(50),
    to_slogic(71),
    to_slogic(63),
    to_slogic(44),
    to_slogic(50),
    to_slogic(50),
    to_slogic(109),
    to_slogic(130),
    to_slogic(115),
    to_slogic(56),
    to_slogic(65),
    to_slogic(76),
    to_slogic(91),
    to_slogic(115),
    to_slogic(117),
    to_slogic(122),
    to_slogic(140),
    to_slogic(122),
    to_slogic(117),
    to_slogic(120),
    to_slogic(141),
    to_slogic(126),
    to_slogic(96),
    to_slogic(96),
    to_slogic(102),
    to_slogic(56),
    to_slogic(68),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(62),
    to_slogic(64),
    to_slogic(56),
    to_slogic(64),
    to_slogic(70),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(62),
    to_slogic(81),
    to_slogic(97),
    to_slogic(109),
    to_slogic(121),
    to_slogic(118),
    to_slogic(124),
    to_slogic(128),
    to_slogic(134),
    to_slogic(142),
    to_slogic(139),
    to_slogic(149),
    to_slogic(146),
    to_slogic(149),
    to_slogic(149),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(165),
    to_slogic(162),
    to_slogic(169),
    to_slogic(165),
    to_slogic(162),
    to_slogic(151),
    to_slogic(149),
    to_slogic(139),
    to_slogic(109),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(75),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(96),
    to_slogic(101),
    to_slogic(75),
    to_slogic(96),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(70),
    to_slogic(69),
    to_slogic(49),
    to_slogic(91),
    to_slogic(176),
    to_slogic(158),
    to_slogic(162),
    to_slogic(143),
    to_slogic(149),
    to_slogic(150),
    to_slogic(156),
    to_slogic(156),
    to_slogic(149),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(156),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(149),
    to_slogic(132),
    to_slogic(144),
    to_slogic(132),
    to_slogic(143),
    to_slogic(130),
    to_slogic(119),
    to_slogic(119),
    to_slogic(143),
    to_slogic(191),
    to_slogic(213),
    to_slogic(223),
    to_slogic(223),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(198),
    to_slogic(197),
    to_slogic(197),
    to_slogic(197),
    to_slogic(183),
    to_slogic(169),
    to_slogic(144),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(75),
    to_slogic(94),
    to_slogic(96),
    to_slogic(117),
    to_slogic(126),
    to_slogic(133),
    to_slogic(144),
    to_slogic(151),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(172),
    to_slogic(157),
    to_slogic(143),
    to_slogic(116),
    to_slogic(81),
    to_slogic(63),
    to_slogic(69),
    to_slogic(92),
    to_slogic(109),
    to_slogic(63),
    to_slogic(56),
    to_slogic(50),
    to_slogic(58),
    to_slogic(89),
    to_slogic(87),
    to_slogic(64),
    to_slogic(56),
    to_slogic(65),
    to_slogic(56),
    to_slogic(71),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(44),
    to_slogic(97),
    to_slogic(140),
    to_slogic(127),
    to_slogic(76),
    to_slogic(65),
    to_slogic(78),
    to_slogic(91),
    to_slogic(109),
    to_slogic(107),
    to_slogic(122),
    to_slogic(132),
    to_slogic(145),
    to_slogic(132),
    to_slogic(117),
    to_slogic(136),
    to_slogic(160),
    to_slogic(107),
    to_slogic(81),
    to_slogic(101),
    to_slogic(89),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(75),
    to_slogic(56),
    to_slogic(42),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(70),
    to_slogic(70),
    to_slogic(49),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(62),
    to_slogic(81),
    to_slogic(97),
    to_slogic(99),
    to_slogic(100),
    to_slogic(109),
    to_slogic(124),
    to_slogic(128),
    to_slogic(119),
    to_slogic(134),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(149),
    to_slogic(151),
    to_slogic(149),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(155),
    to_slogic(149),
    to_slogic(146),
    to_slogic(139),
    to_slogic(102),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(56),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(91),
    to_slogic(96),
    to_slogic(82),
    to_slogic(92),
    to_slogic(82),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(70),
    to_slogic(82),
    to_slogic(49),
    to_slogic(101),
    to_slogic(172),
    to_slogic(155),
    to_slogic(155),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(143),
    to_slogic(150),
    to_slogic(144),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(143),
    to_slogic(133),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(133),
    to_slogic(130),
    to_slogic(119),
    to_slogic(118),
    to_slogic(150),
    to_slogic(198),
    to_slogic(213),
    to_slogic(222),
    to_slogic(223),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(197),
    to_slogic(191),
    to_slogic(176),
    to_slogic(144),
    to_slogic(116),
    to_slogic(94),
    to_slogic(64),
    to_slogic(44),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(92),
    to_slogic(94),
    to_slogic(109),
    to_slogic(117),
    to_slogic(144),
    to_slogic(152),
    to_slogic(155),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(152),
    to_slogic(135),
    to_slogic(109),
    to_slogic(81),
    to_slogic(49),
    to_slogic(81),
    to_slogic(134),
    to_slogic(102),
    to_slogic(102),
    to_slogic(71),
    to_slogic(42),
    to_slogic(68),
    to_slogic(89),
    to_slogic(63),
    to_slogic(68),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(42),
    to_slogic(50),
    to_slogic(42),
    to_slogic(84),
    to_slogic(145),
    to_slogic(140),
    to_slogic(89),
    to_slogic(71),
    to_slogic(84),
    to_slogic(71),
    to_slogic(91),
    to_slogic(120),
    to_slogic(109),
    to_slogic(97),
    to_slogic(130),
    to_slogic(109),
    to_slogic(132),
    to_slogic(140),
    to_slogic(145),
    to_slogic(136),
    to_slogic(136),
    to_slogic(127),
    to_slogic(133),
    to_slogic(68),
    to_slogic(50),
    to_slogic(49),
    to_slogic(50),
    to_slogic(56),
    to_slogic(50),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(64),
    to_slogic(40),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(62),
    to_slogic(75),
    to_slogic(70),
    to_slogic(64),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(63),
    to_slogic(62),
    to_slogic(76),
    to_slogic(89),
    to_slogic(92),
    to_slogic(96),
    to_slogic(119),
    to_slogic(119),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(149),
    to_slogic(151),
    to_slogic(149),
    to_slogic(151),
    to_slogic(161),
    to_slogic(165),
    to_slogic(161),
    to_slogic(152),
    to_slogic(149),
    to_slogic(151),
    to_slogic(149),
    to_slogic(139),
    to_slogic(139),
    to_slogic(130),
    to_slogic(89),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(96),
    to_slogic(101),
    to_slogic(83),
    to_slogic(83),
    to_slogic(82),
    to_slogic(75),
    to_slogic(83),
    to_slogic(92),
    to_slogic(70),
    to_slogic(75),
    to_slogic(56),
    to_slogic(109),
    to_slogic(172),
    to_slogic(150),
    to_slogic(155),
    to_slogic(137),
    to_slogic(124),
    to_slogic(124),
    to_slogic(130),
    to_slogic(137),
    to_slogic(139),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(156),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(133),
    to_slogic(143),
    to_slogic(132),
    to_slogic(119),
    to_slogic(119),
    to_slogic(119),
    to_slogic(166),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(197),
    to_slogic(191),
    to_slogic(183),
    to_slogic(158),
    to_slogic(136),
    to_slogic(94),
    to_slogic(62),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(62),
    to_slogic(94),
    to_slogic(88),
    to_slogic(92),
    to_slogic(116),
    to_slogic(135),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(152),
    to_slogic(135),
    to_slogic(100),
    to_slogic(77),
    to_slogic(89),
    to_slogic(166),
    to_slogic(158),
    to_slogic(88),
    to_slogic(133),
    to_slogic(68),
    to_slogic(42),
    to_slogic(56),
    to_slogic(81),
    to_slogic(63),
    to_slogic(64),
    to_slogic(63),
    to_slogic(56),
    to_slogic(71),
    to_slogic(49),
    to_slogic(56),
    to_slogic(42),
    to_slogic(50),
    to_slogic(44),
    to_slogic(71),
    to_slogic(145),
    to_slogic(145),
    to_slogic(130),
    to_slogic(91),
    to_slogic(91),
    to_slogic(58),
    to_slogic(78),
    to_slogic(120),
    to_slogic(130),
    to_slogic(76),
    to_slogic(109),
    to_slogic(109),
    to_slogic(117),
    to_slogic(155),
    to_slogic(145),
    to_slogic(130),
    to_slogic(126),
    to_slogic(152),
    to_slogic(153),
    to_slogic(115),
    to_slogic(63),
    to_slogic(56),
    to_slogic(50),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(56),
    to_slogic(40),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(64),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(75),
    to_slogic(89),
    to_slogic(62),
    to_slogic(70),
    to_slogic(75),
    to_slogic(92),
    to_slogic(96),
    to_slogic(92),
    to_slogic(101),
    to_slogic(110),
    to_slogic(117),
    to_slogic(119),
    to_slogic(119),
    to_slogic(119),
    to_slogic(127),
    to_slogic(128),
    to_slogic(134),
    to_slogic(142),
    to_slogic(149),
    to_slogic(151),
    to_slogic(151),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(161),
    to_slogic(157),
    to_slogic(157),
    to_slogic(151),
    to_slogic(149),
    to_slogic(139),
    to_slogic(133),
    to_slogic(91),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(96),
    to_slogic(96),
    to_slogic(92),
    to_slogic(83),
    to_slogic(83),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(70),
    to_slogic(77),
    to_slogic(63),
    to_slogic(109),
    to_slogic(176),
    to_slogic(157),
    to_slogic(143),
    to_slogic(118),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(124),
    to_slogic(125),
    to_slogic(130),
    to_slogic(132),
    to_slogic(130),
    to_slogic(132),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(149),
    to_slogic(144),
    to_slogic(143),
    to_slogic(149),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(119),
    to_slogic(119),
    to_slogic(114),
    to_slogic(119),
    to_slogic(171),
    to_slogic(207),
    to_slogic(222),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(205),
    to_slogic(191),
    to_slogic(183),
    to_slogic(161),
    to_slogic(130),
    to_slogic(94),
    to_slogic(64),
    to_slogic(49),
    to_slogic(33),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(40),
    to_slogic(44),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(89),
    to_slogic(82),
    to_slogic(109),
    to_slogic(133),
    to_slogic(144),
    to_slogic(155),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(130),
    to_slogic(109),
    to_slogic(113),
    to_slogic(181),
    to_slogic(158),
    to_slogic(83),
    to_slogic(69),
    to_slogic(143),
    to_slogic(63),
    to_slogic(50),
    to_slogic(49),
    to_slogic(89),
    to_slogic(71),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(50),
    to_slogic(42),
    to_slogic(50),
    to_slogic(71),
    to_slogic(132),
    to_slogic(122),
    to_slogic(145),
    to_slogic(97),
    to_slogic(81),
    to_slogic(71),
    to_slogic(56),
    to_slogic(89),
    to_slogic(113),
    to_slogic(78),
    to_slogic(130),
    to_slogic(140),
    to_slogic(91),
    to_slogic(130),
    to_slogic(155),
    to_slogic(130),
    to_slogic(81),
    to_slogic(75),
    to_slogic(119),
    to_slogic(163),
    to_slogic(127),
    to_slogic(71),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(75),
    to_slogic(64),
    to_slogic(40),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(70),
    to_slogic(81),
    to_slogic(81),
    to_slogic(92),
    to_slogic(102),
    to_slogic(109),
    to_slogic(117),
    to_slogic(126),
    to_slogic(128),
    to_slogic(134),
    to_slogic(133),
    to_slogic(146),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(146),
    to_slogic(134),
    to_slogic(146),
    to_slogic(151),
    to_slogic(151),
    to_slogic(155),
    to_slogic(155),
    to_slogic(151),
    to_slogic(155),
    to_slogic(155),
    to_slogic(162),
    to_slogic(165),
    to_slogic(162),
    to_slogic(172),
    to_slogic(176),
    to_slogic(182),
    to_slogic(185),
    to_slogic(162),
    to_slogic(119),
    to_slogic(95),
    to_slogic(63),
    to_slogic(68),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(96),
    to_slogic(96),
    to_slogic(82),
    to_slogic(96),
    to_slogic(82),
    to_slogic(75),
    to_slogic(88),
    to_slogic(82),
    to_slogic(70),
    to_slogic(69),
    to_slogic(69),
    to_slogic(120),
    to_slogic(165),
    to_slogic(150),
    to_slogic(133),
    to_slogic(107),
    to_slogic(118),
    to_slogic(101),
    to_slogic(107),
    to_slogic(118),
    to_slogic(128),
    to_slogic(118),
    to_slogic(124),
    to_slogic(120),
    to_slogic(125),
    to_slogic(130),
    to_slogic(125),
    to_slogic(132),
    to_slogic(132),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(149),
    to_slogic(133),
    to_slogic(143),
    to_slogic(133),
    to_slogic(130),
    to_slogic(132),
    to_slogic(119),
    to_slogic(114),
    to_slogic(130),
    to_slogic(191),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(205),
    to_slogic(207),
    to_slogic(205),
    to_slogic(197),
    to_slogic(193),
    to_slogic(178),
    to_slogic(158),
    to_slogic(118),
    to_slogic(70),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(62),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(62),
    to_slogic(70),
    to_slogic(75),
    to_slogic(75),
    to_slogic(109),
    to_slogic(130),
    to_slogic(144),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(144),
    to_slogic(134),
    to_slogic(133),
    to_slogic(185),
    to_slogic(158),
    to_slogic(75),
    to_slogic(87),
    to_slogic(68),
    to_slogic(102),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(81),
    to_slogic(81),
    to_slogic(64),
    to_slogic(63),
    to_slogic(75),
    to_slogic(56),
    to_slogic(63),
    to_slogic(75),
    to_slogic(49),
    to_slogic(50),
    to_slogic(44),
    to_slogic(83),
    to_slogic(130),
    to_slogic(122),
    to_slogic(120),
    to_slogic(140),
    to_slogic(89),
    to_slogic(71),
    to_slogic(44),
    to_slogic(58),
    to_slogic(109),
    to_slogic(109),
    to_slogic(145),
    to_slogic(120),
    to_slogic(84),
    to_slogic(109),
    to_slogic(143),
    to_slogic(138),
    to_slogic(115),
    to_slogic(83),
    to_slogic(65),
    to_slogic(149),
    to_slogic(168),
    to_slogic(138),
    to_slogic(71),
    to_slogic(50),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(70),
    to_slogic(82),
    to_slogic(64),
    to_slogic(49),
    to_slogic(40),
    to_slogic(82),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(42),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(70),
    to_slogic(75),
    to_slogic(82),
    to_slogic(102),
    to_slogic(109),
    to_slogic(126),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(134),
    to_slogic(133),
    to_slogic(133),
    to_slogic(133),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(144),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(162),
    to_slogic(165),
    to_slogic(176),
    to_slogic(187),
    to_slogic(193),
    to_slogic(198),
    to_slogic(198),
    to_slogic(189),
    to_slogic(165),
    to_slogic(102),
    to_slogic(68),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(69),
    to_slogic(82),
    to_slogic(101),
    to_slogic(82),
    to_slogic(91),
    to_slogic(83),
    to_slogic(75),
    to_slogic(82),
    to_slogic(92),
    to_slogic(81),
    to_slogic(69),
    to_slogic(69),
    to_slogic(125),
    to_slogic(162),
    to_slogic(157),
    to_slogic(124),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(107),
    to_slogic(107),
    to_slogic(109),
    to_slogic(118),
    to_slogic(119),
    to_slogic(119),
    to_slogic(118),
    to_slogic(118),
    to_slogic(120),
    to_slogic(124),
    to_slogic(125),
    to_slogic(132),
    to_slogic(132),
    to_slogic(139),
    to_slogic(133),
    to_slogic(132),
    to_slogic(144),
    to_slogic(133),
    to_slogic(132),
    to_slogic(132),
    to_slogic(119),
    to_slogic(119),
    to_slogic(118),
    to_slogic(144),
    to_slogic(191),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(205),
    to_slogic(205),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(197),
    to_slogic(183),
    to_slogic(162),
    to_slogic(124),
    to_slogic(82),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(56),
    to_slogic(70),
    to_slogic(75),
    to_slogic(75),
    to_slogic(64),
    to_slogic(63),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(70),
    to_slogic(75),
    to_slogic(75),
    to_slogic(94),
    to_slogic(126),
    to_slogic(143),
    to_slogic(152),
    to_slogic(162),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(182),
    to_slogic(130),
    to_slogic(70),
    to_slogic(75),
    to_slogic(56),
    to_slogic(102),
    to_slogic(89),
    to_slogic(40),
    to_slogic(42),
    to_slogic(42),
    to_slogic(75),
    to_slogic(81),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(95),
    to_slogic(65),
    to_slogic(56),
    to_slogic(56),
    to_slogic(65),
    to_slogic(97),
    to_slogic(122),
    to_slogic(120),
    to_slogic(120),
    to_slogic(130),
    to_slogic(78),
    to_slogic(58),
    to_slogic(84),
    to_slogic(122),
    to_slogic(138),
    to_slogic(140),
    to_slogic(89),
    to_slogic(97),
    to_slogic(97),
    to_slogic(107),
    to_slogic(122),
    to_slogic(102),
    to_slogic(95),
    to_slogic(71),
    to_slogic(110),
    to_slogic(148),
    to_slogic(143),
    to_slogic(138),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(64),
    to_slogic(82),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(68),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(70),
    to_slogic(89),
    to_slogic(92),
    to_slogic(109),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(126),
    to_slogic(124),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(134),
    to_slogic(133),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(146),
    to_slogic(146),
    to_slogic(151),
    to_slogic(165),
    to_slogic(172),
    to_slogic(183),
    to_slogic(182),
    to_slogic(198),
    to_slogic(193),
    to_slogic(198),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(165),
    to_slogic(113),
    to_slogic(81),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(82),
    to_slogic(91),
    to_slogic(109),
    to_slogic(75),
    to_slogic(83),
    to_slogic(83),
    to_slogic(82),
    to_slogic(75),
    to_slogic(83),
    to_slogic(75),
    to_slogic(83),
    to_slogic(69),
    to_slogic(133),
    to_slogic(162),
    to_slogic(143),
    to_slogic(124),
    to_slogic(127),
    to_slogic(124),
    to_slogic(125),
    to_slogic(118),
    to_slogic(119),
    to_slogic(118),
    to_slogic(117),
    to_slogic(109),
    to_slogic(107),
    to_slogic(109),
    to_slogic(107),
    to_slogic(107),
    to_slogic(109),
    to_slogic(118),
    to_slogic(109),
    to_slogic(118),
    to_slogic(124),
    to_slogic(119),
    to_slogic(119),
    to_slogic(125),
    to_slogic(132),
    to_slogic(119),
    to_slogic(132),
    to_slogic(119),
    to_slogic(119),
    to_slogic(119),
    to_slogic(114),
    to_slogic(150),
    to_slogic(197),
    to_slogic(213),
    to_slogic(213),
    to_slogic(205),
    to_slogic(207),
    to_slogic(205),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(205),
    to_slogic(197),
    to_slogic(191),
    to_slogic(183),
    to_slogic(166),
    to_slogic(144),
    to_slogic(88),
    to_slogic(56),
    to_slogic(40),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(70),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(96),
    to_slogic(83),
    to_slogic(75),
    to_slogic(70),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(62),
    to_slogic(62),
    to_slogic(62),
    to_slogic(89),
    to_slogic(121),
    to_slogic(135),
    to_slogic(152),
    to_slogic(157),
    to_slogic(173),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(165),
    to_slogic(165),
    to_slogic(187),
    to_slogic(130),
    to_slogic(76),
    to_slogic(69),
    to_slogic(75),
    to_slogic(75),
    to_slogic(149),
    to_slogic(68),
    to_slogic(40),
    to_slogic(49),
    to_slogic(36),
    to_slogic(63),
    to_slogic(81),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(95),
    to_slogic(88),
    to_slogic(56),
    to_slogic(63),
    to_slogic(58),
    to_slogic(56),
    to_slogic(102),
    to_slogic(130),
    to_slogic(91),
    to_slogic(120),
    to_slogic(122),
    to_slogic(122),
    to_slogic(122),
    to_slogic(140),
    to_slogic(155),
    to_slogic(102),
    to_slogic(78),
    to_slogic(91),
    to_slogic(107),
    to_slogic(91),
    to_slogic(120),
    to_slogic(115),
    to_slogic(76),
    to_slogic(117),
    to_slogic(138),
    to_slogic(143),
    to_slogic(102),
    to_slogic(138),
    to_slogic(127),
    to_slogic(50),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(75),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(82),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(70),
    to_slogic(82),
    to_slogic(92),
    to_slogic(118),
    to_slogic(117),
    to_slogic(124),
    to_slogic(124),
    to_slogic(128),
    to_slogic(117),
    to_slogic(126),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(133),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(144),
    to_slogic(146),
    to_slogic(134),
    to_slogic(146),
    to_slogic(139),
    to_slogic(137),
    to_slogic(149),
    to_slogic(152),
    to_slogic(151),
    to_slogic(173),
    to_slogic(166),
    to_slogic(177),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(198),
    to_slogic(207),
    to_slogic(200),
    to_slogic(198),
    to_slogic(207),
    to_slogic(200),
    to_slogic(170),
    to_slogic(119),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(75),
    to_slogic(83),
    to_slogic(96),
    to_slogic(75),
    to_slogic(83),
    to_slogic(82),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(70),
    to_slogic(75),
    to_slogic(63),
    to_slogic(149),
    to_slogic(150),
    to_slogic(146),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(137),
    to_slogic(130),
    to_slogic(133),
    to_slogic(124),
    to_slogic(118),
    to_slogic(117),
    to_slogic(118),
    to_slogic(107),
    to_slogic(107),
    to_slogic(107),
    to_slogic(107),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(107),
    to_slogic(107),
    to_slogic(118),
    to_slogic(107),
    to_slogic(102),
    to_slogic(118),
    to_slogic(118),
    to_slogic(118),
    to_slogic(118),
    to_slogic(109),
    to_slogic(109),
    to_slogic(143),
    to_slogic(197),
    to_slogic(207),
    to_slogic(213),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(197),
    to_slogic(183),
    to_slogic(172),
    to_slogic(130),
    to_slogic(82),
    to_slogic(56),
    to_slogic(44),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(70),
    to_slogic(89),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(126),
    to_slogic(119),
    to_slogic(102),
    to_slogic(83),
    to_slogic(82),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(76),
    to_slogic(100),
    to_slogic(130),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(179),
    to_slogic(187),
    to_slogic(173),
    to_slogic(144),
    to_slogic(116),
    to_slogic(82),
    to_slogic(69),
    to_slogic(101),
    to_slogic(143),
    to_slogic(96),
    to_slogic(49),
    to_slogic(42),
    to_slogic(40),
    to_slogic(42),
    to_slogic(49),
    to_slogic(63),
    to_slogic(81),
    to_slogic(75),
    to_slogic(49),
    to_slogic(42),
    to_slogic(50),
    to_slogic(83),
    to_slogic(102),
    to_slogic(75),
    to_slogic(65),
    to_slogic(83),
    to_slogic(42),
    to_slogic(56),
    to_slogic(130),
    to_slogic(120),
    to_slogic(89),
    to_slogic(71),
    to_slogic(89),
    to_slogic(97),
    to_slogic(143),
    to_slogic(120),
    to_slogic(78),
    to_slogic(91),
    to_slogic(97),
    to_slogic(91),
    to_slogic(122),
    to_slogic(109),
    to_slogic(107),
    to_slogic(107),
    to_slogic(115),
    to_slogic(166),
    to_slogic(133),
    to_slogic(89),
    to_slogic(75),
    to_slogic(143),
    to_slogic(81),
    to_slogic(42),
    to_slogic(56),
    to_slogic(63),
    to_slogic(82),
    to_slogic(56),
    to_slogic(42),
    to_slogic(56),
    to_slogic(82),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(92),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(128),
    to_slogic(126),
    to_slogic(126),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(133),
    to_slogic(142),
    to_slogic(144),
    to_slogic(146),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(144),
    to_slogic(152),
    to_slogic(151),
    to_slogic(173),
    to_slogic(172),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(198),
    to_slogic(198),
    to_slogic(198),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(207),
    to_slogic(200),
    to_slogic(177),
    to_slogic(114),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(49),
    to_slogic(75),
    to_slogic(75),
    to_slogic(96),
    to_slogic(75),
    to_slogic(83),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(70),
    to_slogic(69),
    to_slogic(149),
    to_slogic(152),
    to_slogic(143),
    to_slogic(130),
    to_slogic(139),
    to_slogic(130),
    to_slogic(130),
    to_slogic(143),
    to_slogic(130),
    to_slogic(125),
    to_slogic(124),
    to_slogic(125),
    to_slogic(127),
    to_slogic(118),
    to_slogic(119),
    to_slogic(107),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(101),
    to_slogic(107),
    to_slogic(107),
    to_slogic(102),
    to_slogic(96),
    to_slogic(91),
    to_slogic(137),
    to_slogic(191),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(191),
    to_slogic(166),
    to_slogic(130),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(70),
    to_slogic(70),
    to_slogic(75),
    to_slogic(89),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(133),
    to_slogic(133),
    to_slogic(119),
    to_slogic(102),
    to_slogic(91),
    to_slogic(82),
    to_slogic(75),
    to_slogic(64),
    to_slogic(70),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(70),
    to_slogic(100),
    to_slogic(130),
    to_slogic(144),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(173),
    to_slogic(157),
    to_slogic(139),
    to_slogic(109),
    to_slogic(82),
    to_slogic(102),
    to_slogic(125),
    to_slogic(158),
    to_slogic(56),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(50),
    to_slogic(81),
    to_slogic(107),
    to_slogic(40),
    to_slogic(36),
    to_slogic(50),
    to_slogic(81),
    to_slogic(107),
    to_slogic(75),
    to_slogic(81),
    to_slogic(89),
    to_slogic(42),
    to_slogic(42),
    to_slogic(71),
    to_slogic(130),
    to_slogic(130),
    to_slogic(109),
    to_slogic(91),
    to_slogic(89),
    to_slogic(127),
    to_slogic(76),
    to_slogic(84),
    to_slogic(109),
    to_slogic(107),
    to_slogic(107),
    to_slogic(97),
    to_slogic(130),
    to_slogic(117),
    to_slogic(115),
    to_slogic(120),
    to_slogic(134),
    to_slogic(138),
    to_slogic(89),
    to_slogic(65),
    to_slogic(89),
    to_slogic(143),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(75),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(75),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(75),
    to_slogic(94),
    to_slogic(102),
    to_slogic(116),
    to_slogic(116),
    to_slogic(124),
    to_slogic(117),
    to_slogic(124),
    to_slogic(128),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(133),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(139),
    to_slogic(146),
    to_slogic(144),
    to_slogic(149),
    to_slogic(151),
    to_slogic(157),
    to_slogic(172),
    to_slogic(177),
    to_slogic(183),
    to_slogic(193),
    to_slogic(191),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(198),
    to_slogic(207),
    to_slogic(198),
    to_slogic(207),
    to_slogic(200),
    to_slogic(204),
    to_slogic(207),
    to_slogic(204),
    to_slogic(153),
    to_slogic(81),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(69),
    to_slogic(82),
    to_slogic(96),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(70),
    to_slogic(75),
    to_slogic(70),
    to_slogic(69),
    to_slogic(69),
    to_slogic(69),
    to_slogic(149),
    to_slogic(152),
    to_slogic(139),
    to_slogic(141),
    to_slogic(143),
    to_slogic(139),
    to_slogic(143),
    to_slogic(139),
    to_slogic(143),
    to_slogic(137),
    to_slogic(139),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(120),
    to_slogic(118),
    to_slogic(117),
    to_slogic(109),
    to_slogic(107),
    to_slogic(101),
    to_slogic(96),
    to_slogic(96),
    to_slogic(101),
    to_slogic(91),
    to_slogic(91),
    to_slogic(96),
    to_slogic(107),
    to_slogic(118),
    to_slogic(101),
    to_slogic(82),
    to_slogic(75),
    to_slogic(124),
    to_slogic(191),
    to_slogic(205),
    to_slogic(207),
    to_slogic(205),
    to_slogic(205),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(197),
    to_slogic(191),
    to_slogic(172),
    to_slogic(136),
    to_slogic(75),
    to_slogic(40),
    to_slogic(49),
    to_slogic(70),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(82),
    to_slogic(143),
    to_slogic(143),
    to_slogic(133),
    to_slogic(133),
    to_slogic(114),
    to_slogic(101),
    to_slogic(83),
    to_slogic(82),
    to_slogic(75),
    to_slogic(70),
    to_slogic(49),
    to_slogic(44),
    to_slogic(70),
    to_slogic(100),
    to_slogic(126),
    to_slogic(151),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(152),
    to_slogic(143),
    to_slogic(117),
    to_slogic(110),
    to_slogic(126),
    to_slogic(144),
    to_slogic(109),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(42),
    to_slogic(42),
    to_slogic(71),
    to_slogic(81),
    to_slogic(107),
    to_slogic(42),
    to_slogic(36),
    to_slogic(50),
    to_slogic(95),
    to_slogic(126),
    to_slogic(71),
    to_slogic(97),
    to_slogic(81),
    to_slogic(49),
    to_slogic(42),
    to_slogic(71),
    to_slogic(89),
    to_slogic(89),
    to_slogic(120),
    to_slogic(107),
    to_slogic(130),
    to_slogic(120),
    to_slogic(71),
    to_slogic(78),
    to_slogic(95),
    to_slogic(117),
    to_slogic(115),
    to_slogic(97),
    to_slogic(115),
    to_slogic(145),
    to_slogic(122),
    to_slogic(130),
    to_slogic(114),
    to_slogic(133),
    to_slogic(127),
    to_slogic(56),
    to_slogic(83),
    to_slogic(119),
    to_slogic(107),
    to_slogic(56),
    to_slogic(63),
    to_slogic(64),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(82),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(70),
    to_slogic(69),
    to_slogic(62),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(96),
    to_slogic(102),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(128),
    to_slogic(126),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(146),
    to_slogic(146),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(177),
    to_slogic(187),
    to_slogic(187),
    to_slogic(193),
    to_slogic(183),
    to_slogic(193),
    to_slogic(191),
    to_slogic(193),
    to_slogic(198),
    to_slogic(198),
    to_slogic(198),
    to_slogic(207),
    to_slogic(200),
    to_slogic(207),
    to_slogic(204),
    to_slogic(211),
    to_slogic(185),
    to_slogic(102),
    to_slogic(49),
    to_slogic(40),
    to_slogic(64),
    to_slogic(64),
    to_slogic(96),
    to_slogic(69),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(64),
    to_slogic(75),
    to_slogic(155),
    to_slogic(155),
    to_slogic(137),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(133),
    to_slogic(139),
    to_slogic(132),
    to_slogic(139),
    to_slogic(132),
    to_slogic(125),
    to_slogic(125),
    to_slogic(118),
    to_slogic(119),
    to_slogic(107),
    to_slogic(107),
    to_slogic(101),
    to_slogic(96),
    to_slogic(91),
    to_slogic(94),
    to_slogic(107),
    to_slogic(124),
    to_slogic(118),
    to_slogic(118),
    to_slogic(88),
    to_slogic(75),
    to_slogic(118),
    to_slogic(191),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(183),
    to_slogic(161),
    to_slogic(118),
    to_slogic(75),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(94),
    to_slogic(82),
    to_slogic(92),
    to_slogic(82),
    to_slogic(127),
    to_slogic(133),
    to_slogic(149),
    to_slogic(127),
    to_slogic(133),
    to_slogic(119),
    to_slogic(109),
    to_slogic(96),
    to_slogic(88),
    to_slogic(75),
    to_slogic(49),
    to_slogic(44),
    to_slogic(70),
    to_slogic(100),
    to_slogic(130),
    to_slogic(146),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(165),
    to_slogic(152),
    to_slogic(139),
    to_slogic(133),
    to_slogic(155),
    to_slogic(126),
    to_slogic(120),
    to_slogic(68),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(36),
    to_slogic(42),
    to_slogic(81),
    to_slogic(115),
    to_slogic(120),
    to_slogic(91),
    to_slogic(78),
    to_slogic(97),
    to_slogic(120),
    to_slogic(83),
    to_slogic(71),
    to_slogic(75),
    to_slogic(71),
    to_slogic(44),
    to_slogic(58),
    to_slogic(107),
    to_slogic(71),
    to_slogic(58),
    to_slogic(97),
    to_slogic(120),
    to_slogic(95),
    to_slogic(71),
    to_slogic(71),
    to_slogic(78),
    to_slogic(76),
    to_slogic(102),
    to_slogic(122),
    to_slogic(115),
    to_slogic(122),
    to_slogic(145),
    to_slogic(140),
    to_slogic(127),
    to_slogic(107),
    to_slogic(68),
    to_slogic(119),
    to_slogic(102),
    to_slogic(50),
    to_slogic(83),
    to_slogic(143),
    to_slogic(71),
    to_slogic(56),
    to_slogic(64),
    to_slogic(50),
    to_slogic(49),
    to_slogic(49),
    to_slogic(82),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(64),
    to_slogic(82),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(75),
    to_slogic(96),
    to_slogic(101),
    to_slogic(115),
    to_slogic(115),
    to_slogic(117),
    to_slogic(124),
    to_slogic(128),
    to_slogic(124),
    to_slogic(128),
    to_slogic(128),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(146),
    to_slogic(144),
    to_slogic(139),
    to_slogic(134),
    to_slogic(134),
    to_slogic(146),
    to_slogic(146),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(187),
    to_slogic(183),
    to_slogic(193),
    to_slogic(183),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(193),
    to_slogic(198),
    to_slogic(207),
    to_slogic(198),
    to_slogic(207),
    to_slogic(204),
    to_slogic(207),
    to_slogic(211),
    to_slogic(213),
    to_slogic(196),
    to_slogic(119),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(91),
    to_slogic(64),
    to_slogic(68),
    to_slogic(70),
    to_slogic(64),
    to_slogic(75),
    to_slogic(70),
    to_slogic(70),
    to_slogic(56),
    to_slogic(83),
    to_slogic(162),
    to_slogic(143),
    to_slogic(137),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(133),
    to_slogic(139),
    to_slogic(132),
    to_slogic(130),
    to_slogic(125),
    to_slogic(124),
    to_slogic(125),
    to_slogic(118),
    to_slogic(118),
    to_slogic(109),
    to_slogic(107),
    to_slogic(101),
    to_slogic(101),
    to_slogic(102),
    to_slogic(118),
    to_slogic(136),
    to_slogic(116),
    to_slogic(88),
    to_slogic(82),
    to_slogic(144),
    to_slogic(197),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(197),
    to_slogic(172),
    to_slogic(107),
    to_slogic(63),
    to_slogic(44),
    to_slogic(49),
    to_slogic(75),
    to_slogic(82),
    to_slogic(89),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(94),
    to_slogic(92),
    to_slogic(82),
    to_slogic(81),
    to_slogic(82),
    to_slogic(133),
    to_slogic(133),
    to_slogic(153),
    to_slogic(153),
    to_slogic(149),
    to_slogic(133),
    to_slogic(119),
    to_slogic(114),
    to_slogic(96),
    to_slogic(75),
    to_slogic(56),
    to_slogic(44),
    to_slogic(62),
    to_slogic(100),
    to_slogic(128),
    to_slogic(144),
    to_slogic(162),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(173),
    to_slogic(165),
    to_slogic(152),
    to_slogic(139),
    to_slogic(169),
    to_slogic(185),
    to_slogic(101),
    to_slogic(101),
    to_slogic(69),
    to_slogic(50),
    to_slogic(40),
    to_slogic(42),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(56),
    to_slogic(71),
    to_slogic(81),
    to_slogic(95),
    to_slogic(113),
    to_slogic(121),
    to_slogic(75),
    to_slogic(75),
    to_slogic(71),
    to_slogic(65),
    to_slogic(71),
    to_slogic(76),
    to_slogic(113),
    to_slogic(89),
    to_slogic(50),
    to_slogic(58),
    to_slogic(120),
    to_slogic(81),
    to_slogic(71),
    to_slogic(65),
    to_slogic(58),
    to_slogic(83),
    to_slogic(91),
    to_slogic(84),
    to_slogic(107),
    to_slogic(122),
    to_slogic(130),
    to_slogic(140),
    to_slogic(140),
    to_slogic(140),
    to_slogic(138),
    to_slogic(56),
    to_slogic(56),
    to_slogic(152),
    to_slogic(89),
    to_slogic(56),
    to_slogic(114),
    to_slogic(119),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(82),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(70),
    to_slogic(92),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(82),
    to_slogic(82),
    to_slogic(109),
    to_slogic(117),
    to_slogic(117),
    to_slogic(124),
    to_slogic(126),
    to_slogic(126),
    to_slogic(117),
    to_slogic(128),
    to_slogic(128),
    to_slogic(133),
    to_slogic(139),
    to_slogic(142),
    to_slogic(144),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(151),
    to_slogic(157),
    to_slogic(162),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(177),
    to_slogic(187),
    to_slogic(187),
    to_slogic(183),
    to_slogic(193),
    to_slogic(191),
    to_slogic(187),
    to_slogic(193),
    to_slogic(198),
    to_slogic(198),
    to_slogic(198),
    to_slogic(207),
    to_slogic(200),
    to_slogic(207),
    to_slogic(211),
    to_slogic(207),
    to_slogic(214),
    to_slogic(204),
    to_slogic(133),
    to_slogic(56),
    to_slogic(49),
    to_slogic(82),
    to_slogic(56),
    to_slogic(64),
    to_slogic(64),
    to_slogic(64),
    to_slogic(75),
    to_slogic(70),
    to_slogic(64),
    to_slogic(46),
    to_slogic(83),
    to_slogic(155),
    to_slogic(152),
    to_slogic(139),
    to_slogic(150),
    to_slogic(144),
    to_slogic(150),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(132),
    to_slogic(132),
    to_slogic(139),
    to_slogic(132),
    to_slogic(132),
    to_slogic(125),
    to_slogic(125),
    to_slogic(120),
    to_slogic(118),
    to_slogic(120),
    to_slogic(109),
    to_slogic(102),
    to_slogic(118),
    to_slogic(130),
    to_slogic(136),
    to_slogic(102),
    to_slogic(94),
    to_slogic(102),
    to_slogic(158),
    to_slogic(205),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(205),
    to_slogic(197),
    to_slogic(191),
    to_slogic(136),
    to_slogic(75),
    to_slogic(40),
    to_slogic(56),
    to_slogic(75),
    to_slogic(88),
    to_slogic(92),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(94),
    to_slogic(96),
    to_slogic(94),
    to_slogic(96),
    to_slogic(88),
    to_slogic(82),
    to_slogic(92),
    to_slogic(133),
    to_slogic(127),
    to_slogic(149),
    to_slogic(143),
    to_slogic(153),
    to_slogic(149),
    to_slogic(143),
    to_slogic(119),
    to_slogic(102),
    to_slogic(82),
    to_slogic(64),
    to_slogic(44),
    to_slogic(62),
    to_slogic(100),
    to_slogic(126),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(165),
    to_slogic(144),
    to_slogic(146),
    to_slogic(200),
    to_slogic(176),
    to_slogic(101),
    to_slogic(81),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(50),
    to_slogic(63),
    to_slogic(63),
    to_slogic(42),
    to_slogic(56),
    to_slogic(81),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(71),
    to_slogic(89),
    to_slogic(95),
    to_slogic(81),
    to_slogic(50),
    to_slogic(42),
    to_slogic(89),
    to_slogic(138),
    to_slogic(50),
    to_slogic(65),
    to_slogic(76),
    to_slogic(65),
    to_slogic(65),
    to_slogic(97),
    to_slogic(97),
    to_slogic(91),
    to_slogic(107),
    to_slogic(122),
    to_slogic(138),
    to_slogic(130),
    to_slogic(153),
    to_slogic(152),
    to_slogic(97),
    to_slogic(44),
    to_slogic(114),
    to_slogic(162),
    to_slogic(71),
    to_slogic(95),
    to_slogic(148),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(49),
    to_slogic(82),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(70),
    to_slogic(75),
    to_slogic(89),
    to_slogic(92),
    to_slogic(49),
    to_slogic(44),
    to_slogic(70),
    to_slogic(82),
    to_slogic(117),
    to_slogic(115),
    to_slogic(121),
    to_slogic(130),
    to_slogic(117),
    to_slogic(118),
    to_slogic(119),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(133),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(139),
    to_slogic(139),
    to_slogic(142),
    to_slogic(146),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(177),
    to_slogic(176),
    to_slogic(177),
    to_slogic(183),
    to_slogic(187),
    to_slogic(183),
    to_slogic(193),
    to_slogic(193),
    to_slogic(197),
    to_slogic(193),
    to_slogic(198),
    to_slogic(198),
    to_slogic(207),
    to_slogic(200),
    to_slogic(207),
    to_slogic(211),
    to_slogic(213),
    to_slogic(213),
    to_slogic(204),
    to_slogic(119),
    to_slogic(56),
    to_slogic(75),
    to_slogic(64),
    to_slogic(62),
    to_slogic(56),
    to_slogic(75),
    to_slogic(82),
    to_slogic(69),
    to_slogic(70),
    to_slogic(49),
    to_slogic(91),
    to_slogic(162),
    to_slogic(143),
    to_slogic(132),
    to_slogic(149),
    to_slogic(150),
    to_slogic(149),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(132),
    to_slogic(144),
    to_slogic(143),
    to_slogic(133),
    to_slogic(143),
    to_slogic(132),
    to_slogic(125),
    to_slogic(132),
    to_slogic(125),
    to_slogic(119),
    to_slogic(119),
    to_slogic(114),
    to_slogic(118),
    to_slogic(118),
    to_slogic(130),
    to_slogic(136),
    to_slogic(116),
    to_slogic(109),
    to_slogic(118),
    to_slogic(183),
    to_slogic(207),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(205),
    to_slogic(196),
    to_slogic(176),
    to_slogic(118),
    to_slogic(49),
    to_slogic(49),
    to_slogic(70),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(82),
    to_slogic(82),
    to_slogic(92),
    to_slogic(96),
    to_slogic(109),
    to_slogic(101),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(119),
    to_slogic(126),
    to_slogic(133),
    to_slogic(153),
    to_slogic(153),
    to_slogic(153),
    to_slogic(149),
    to_slogic(133),
    to_slogic(132),
    to_slogic(96),
    to_slogic(64),
    to_slogic(44),
    to_slogic(70),
    to_slogic(99),
    to_slogic(126),
    to_slogic(152),
    to_slogic(162),
    to_slogic(173),
    to_slogic(173),
    to_slogic(176),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(172),
    to_slogic(165),
    to_slogic(152),
    to_slogic(146),
    to_slogic(200),
    to_slogic(152),
    to_slogic(126),
    to_slogic(133),
    to_slogic(42),
    to_slogic(40),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(68),
    to_slogic(68),
    to_slogic(49),
    to_slogic(63),
    to_slogic(68),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(65),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(89),
    to_slogic(120),
    to_slogic(71),
    to_slogic(44),
    to_slogic(71),
    to_slogic(76),
    to_slogic(76),
    to_slogic(76),
    to_slogic(107),
    to_slogic(97),
    to_slogic(89),
    to_slogic(115),
    to_slogic(140),
    to_slogic(130),
    to_slogic(138),
    to_slogic(120),
    to_slogic(127),
    to_slogic(84),
    to_slogic(89),
    to_slogic(162),
    to_slogic(127),
    to_slogic(81),
    to_slogic(119),
    to_slogic(95),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(50),
    to_slogic(56),
    to_slogic(64),
    to_slogic(68),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(64),
    to_slogic(83),
    to_slogic(64),
    to_slogic(75),
    to_slogic(109),
    to_slogic(96),
    to_slogic(64),
    to_slogic(49),
    to_slogic(70),
    to_slogic(83),
    to_slogic(119),
    to_slogic(117),
    to_slogic(118),
    to_slogic(117),
    to_slogic(117),
    to_slogic(117),
    to_slogic(134),
    to_slogic(134),
    to_slogic(133),
    to_slogic(139),
    to_slogic(133),
    to_slogic(142),
    to_slogic(144),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(151),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(176),
    to_slogic(177),
    to_slogic(183),
    to_slogic(183),
    to_slogic(187),
    to_slogic(191),
    to_slogic(193),
    to_slogic(193),
    to_slogic(205),
    to_slogic(198),
    to_slogic(198),
    to_slogic(207),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(204),
    to_slogic(109),
    to_slogic(56),
    to_slogic(62),
    to_slogic(49),
    to_slogic(56),
    to_slogic(70),
    to_slogic(64),
    to_slogic(75),
    to_slogic(69),
    to_slogic(46),
    to_slogic(109),
    to_slogic(157),
    to_slogic(143),
    to_slogic(137),
    to_slogic(144),
    to_slogic(149),
    to_slogic(150),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(132),
    to_slogic(132),
    to_slogic(141),
    to_slogic(132),
    to_slogic(139),
    to_slogic(132),
    to_slogic(132),
    to_slogic(125),
    to_slogic(132),
    to_slogic(125),
    to_slogic(119),
    to_slogic(118),
    to_slogic(118),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(102),
    to_slogic(144),
    to_slogic(191),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(205),
    to_slogic(183),
    to_slogic(144),
    to_slogic(94),
    to_slogic(56),
    to_slogic(63),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(92),
    to_slogic(92),
    to_slogic(101),
    to_slogic(107),
    to_slogic(107),
    to_slogic(102),
    to_slogic(96),
    to_slogic(82),
    to_slogic(92),
    to_slogic(96),
    to_slogic(91),
    to_slogic(102),
    to_slogic(133),
    to_slogic(143),
    to_slogic(153),
    to_slogic(153),
    to_slogic(153),
    to_slogic(153),
    to_slogic(133),
    to_slogic(102),
    to_slogic(70),
    to_slogic(44),
    to_slogic(62),
    to_slogic(94),
    to_slogic(130),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(172),
    to_slogic(152),
    to_slogic(144),
    to_slogic(176),
    to_slogic(126),
    to_slogic(83),
    to_slogic(102),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(68),
    to_slogic(64),
    to_slogic(63),
    to_slogic(49),
    to_slogic(50),
    to_slogic(42),
    to_slogic(56),
    to_slogic(96),
    to_slogic(68),
    to_slogic(56),
    to_slogic(40),
    to_slogic(42),
    to_slogic(49),
    to_slogic(81),
    to_slogic(42),
    to_slogic(44),
    to_slogic(81),
    to_slogic(102),
    to_slogic(65),
    to_slogic(56),
    to_slogic(65),
    to_slogic(76),
    to_slogic(76),
    to_slogic(89),
    to_slogic(109),
    to_slogic(91),
    to_slogic(102),
    to_slogic(140),
    to_slogic(136),
    to_slogic(130),
    to_slogic(115),
    to_slogic(136),
    to_slogic(115),
    to_slogic(102),
    to_slogic(95),
    to_slogic(138),
    to_slogic(83),
    to_slogic(91),
    to_slogic(152),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(82),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(64),
    to_slogic(82),
    to_slogic(109),
    to_slogic(100),
    to_slogic(70),
    to_slogic(44),
    to_slogic(56),
    to_slogic(82),
    to_slogic(119),
    to_slogic(124),
    to_slogic(109),
    to_slogic(116),
    to_slogic(128),
    to_slogic(134),
    to_slogic(128),
    to_slogic(134),
    to_slogic(139),
    to_slogic(142),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(177),
    to_slogic(178),
    to_slogic(177),
    to_slogic(177),
    to_slogic(177),
    to_slogic(183),
    to_slogic(187),
    to_slogic(191),
    to_slogic(193),
    to_slogic(198),
    to_slogic(198),
    to_slogic(207),
    to_slogic(200),
    to_slogic(207),
    to_slogic(211),
    to_slogic(204),
    to_slogic(214),
    to_slogic(214),
    to_slogic(213),
    to_slogic(196),
    to_slogic(87),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(64),
    to_slogic(62),
    to_slogic(63),
    to_slogic(63),
    to_slogic(49),
    to_slogic(118),
    to_slogic(150),
    to_slogic(137),
    to_slogic(143),
    to_slogic(149),
    to_slogic(150),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(132),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(133),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(119),
    to_slogic(125),
    to_slogic(125),
    to_slogic(124),
    to_slogic(124),
    to_slogic(136),
    to_slogic(136),
    to_slogic(130),
    to_slogic(118),
    to_slogic(158),
    to_slogic(197),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(191),
    to_slogic(169),
    to_slogic(126),
    to_slogic(82),
    to_slogic(63),
    to_slogic(82),
    to_slogic(100),
    to_slogic(83),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(101),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(94),
    to_slogic(96),
    to_slogic(92),
    to_slogic(102),
    to_slogic(101),
    to_slogic(56),
    to_slogic(81),
    to_slogic(114),
    to_slogic(133),
    to_slogic(143),
    to_slogic(165),
    to_slogic(165),
    to_slogic(153),
    to_slogic(149),
    to_slogic(119),
    to_slogic(75),
    to_slogic(40),
    to_slogic(62),
    to_slogic(99),
    to_slogic(126),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(152),
    to_slogic(144),
    to_slogic(176),
    to_slogic(120),
    to_slogic(87),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(68),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(71),
    to_slogic(102),
    to_slogic(71),
    to_slogic(71),
    to_slogic(56),
    to_slogic(42),
    to_slogic(42),
    to_slogic(95),
    to_slogic(56),
    to_slogic(42),
    to_slogic(71),
    to_slogic(97),
    to_slogic(89),
    to_slogic(56),
    to_slogic(71),
    to_slogic(76),
    to_slogic(71),
    to_slogic(78),
    to_slogic(102),
    to_slogic(97),
    to_slogic(107),
    to_slogic(130),
    to_slogic(120),
    to_slogic(130),
    to_slogic(136),
    to_slogic(145),
    to_slogic(138),
    to_slogic(121),
    to_slogic(63),
    to_slogic(119),
    to_slogic(138),
    to_slogic(68),
    to_slogic(181),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(75),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(75),
    to_slogic(64),
    to_slogic(92),
    to_slogic(116),
    to_slogic(116),
    to_slogic(89),
    to_slogic(44),
    to_slogic(56),
    to_slogic(82),
    to_slogic(109),
    to_slogic(109),
    to_slogic(118),
    to_slogic(126),
    to_slogic(139),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(142),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(177),
    to_slogic(177),
    to_slogic(183),
    to_slogic(183),
    to_slogic(183),
    to_slogic(187),
    to_slogic(193),
    to_slogic(197),
    to_slogic(198),
    to_slogic(198),
    to_slogic(207),
    to_slogic(200),
    to_slogic(207),
    to_slogic(211),
    to_slogic(213),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(165),
    to_slogic(69),
    to_slogic(40),
    to_slogic(44),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(46),
    to_slogic(137),
    to_slogic(152),
    to_slogic(137),
    to_slogic(143),
    to_slogic(143),
    to_slogic(150),
    to_slogic(150),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(133),
    to_slogic(143),
    to_slogic(133),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(119),
    to_slogic(125),
    to_slogic(136),
    to_slogic(136),
    to_slogic(136),
    to_slogic(130),
    to_slogic(130),
    to_slogic(176),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(205),
    to_slogic(191),
    to_slogic(144),
    to_slogic(102),
    to_slogic(69),
    to_slogic(75),
    to_slogic(83),
    to_slogic(96),
    to_slogic(92),
    to_slogic(92),
    to_slogic(94),
    to_slogic(96),
    to_slogic(101),
    to_slogic(107),
    to_slogic(107),
    to_slogic(102),
    to_slogic(96),
    to_slogic(92),
    to_slogic(96),
    to_slogic(96),
    to_slogic(101),
    to_slogic(40),
    to_slogic(63),
    to_slogic(95),
    to_slogic(119),
    to_slogic(153),
    to_slogic(162),
    to_slogic(162),
    to_slogic(165),
    to_slogic(158),
    to_slogic(119),
    to_slogic(88),
    to_slogic(44),
    to_slogic(62),
    to_slogic(94),
    to_slogic(134),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(172),
    to_slogic(152),
    to_slogic(144),
    to_slogic(187),
    to_slogic(121),
    to_slogic(83),
    to_slogic(71),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(42),
    to_slogic(89),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(42),
    to_slogic(42),
    to_slogic(81),
    to_slogic(107),
    to_slogic(56),
    to_slogic(68),
    to_slogic(63),
    to_slogic(40),
    to_slogic(42),
    to_slogic(81),
    to_slogic(89),
    to_slogic(44),
    to_slogic(56),
    to_slogic(89),
    to_slogic(71),
    to_slogic(91),
    to_slogic(58),
    to_slogic(84),
    to_slogic(89),
    to_slogic(76),
    to_slogic(76),
    to_slogic(97),
    to_slogic(107),
    to_slogic(102),
    to_slogic(107),
    to_slogic(122),
    to_slogic(130),
    to_slogic(153),
    to_slogic(163),
    to_slogic(121),
    to_slogic(50),
    to_slogic(49),
    to_slogic(143),
    to_slogic(83),
    to_slogic(196),
    to_slogic(68),
    to_slogic(33),
    to_slogic(40),
    to_slogic(40),
    to_slogic(64),
    to_slogic(64),
    to_slogic(62),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(64),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(63),
    to_slogic(62),
    to_slogic(99),
    to_slogic(116),
    to_slogic(116),
    to_slogic(89),
    to_slogic(44),
    to_slogic(56),
    to_slogic(75),
    to_slogic(102),
    to_slogic(118),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(162),
    to_slogic(162),
    to_slogic(172),
    to_slogic(173),
    to_slogic(172),
    to_slogic(177),
    to_slogic(178),
    to_slogic(187),
    to_slogic(183),
    to_slogic(193),
    to_slogic(187),
    to_slogic(197),
    to_slogic(193),
    to_slogic(198),
    to_slogic(207),
    to_slogic(200),
    to_slogic(204),
    to_slogic(207),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(213),
    to_slogic(132),
    to_slogic(40),
    to_slogic(44),
    to_slogic(62),
    to_slogic(44),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(139),
    to_slogic(143),
    to_slogic(137),
    to_slogic(143),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(139),
    to_slogic(144),
    to_slogic(132),
    to_slogic(133),
    to_slogic(132),
    to_slogic(125),
    to_slogic(125),
    to_slogic(130),
    to_slogic(124),
    to_slogic(130),
    to_slogic(136),
    to_slogic(136),
    to_slogic(136),
    to_slogic(136),
    to_slogic(183),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(205),
    to_slogic(176),
    to_slogic(130),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(96),
    to_slogic(92),
    to_slogic(96),
    to_slogic(96),
    to_slogic(96),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(102),
    to_slogic(92),
    to_slogic(96),
    to_slogic(92),
    to_slogic(101),
    to_slogic(109),
    to_slogic(101),
    to_slogic(33),
    to_slogic(49),
    to_slogic(83),
    to_slogic(114),
    to_slogic(153),
    to_slogic(162),
    to_slogic(170),
    to_slogic(170),
    to_slogic(153),
    to_slogic(132),
    to_slogic(96),
    to_slogic(49),
    to_slogic(49),
    to_slogic(89),
    to_slogic(130),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(165),
    to_slogic(156),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(102),
    to_slogic(83),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(68),
    to_slogic(68),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(75),
    to_slogic(120),
    to_slogic(56),
    to_slogic(63),
    to_slogic(68),
    to_slogic(40),
    to_slogic(36),
    to_slogic(50),
    to_slogic(81),
    to_slogic(71),
    to_slogic(42),
    to_slogic(89),
    to_slogic(58),
    to_slogic(89),
    to_slogic(91),
    to_slogic(78),
    to_slogic(102),
    to_slogic(97),
    to_slogic(78),
    to_slogic(76),
    to_slogic(102),
    to_slogic(97),
    to_slogic(115),
    to_slogic(130),
    to_slogic(115),
    to_slogic(140),
    to_slogic(168),
    to_slogic(119),
    to_slogic(56),
    to_slogic(42),
    to_slogic(83),
    to_slogic(107),
    to_slogic(197),
    to_slogic(89),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(75),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(68),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(62),
    to_slogic(70),
    to_slogic(109),
    to_slogic(116),
    to_slogic(109),
    to_slogic(89),
    to_slogic(44),
    to_slogic(49),
    to_slogic(82),
    to_slogic(101),
    to_slogic(121),
    to_slogic(124),
    to_slogic(126),
    to_slogic(134),
    to_slogic(134),
    to_slogic(134),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(146),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(178),
    to_slogic(177),
    to_slogic(177),
    to_slogic(187),
    to_slogic(183),
    to_slogic(193),
    to_slogic(191),
    to_slogic(193),
    to_slogic(198),
    to_slogic(198),
    to_slogic(198),
    to_slogic(207),
    to_slogic(207),
    to_slogic(204),
    to_slogic(211),
    to_slogic(213),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(200),
    to_slogic(69),
    to_slogic(40),
    to_slogic(62),
    to_slogic(44),
    to_slogic(56),
    to_slogic(33),
    to_slogic(63),
    to_slogic(143),
    to_slogic(144),
    to_slogic(130),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(143),
    to_slogic(133),
    to_slogic(132),
    to_slogic(144),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(125),
    to_slogic(124),
    to_slogic(130),
    to_slogic(136),
    to_slogic(156),
    to_slogic(161),
    to_slogic(172),
    to_slogic(191),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(207),
    to_slogic(203),
    to_slogic(161),
    to_slogic(102),
    to_slogic(75),
    to_slogic(82),
    to_slogic(92),
    to_slogic(94),
    to_slogic(92),
    to_slogic(96),
    to_slogic(109),
    to_slogic(101),
    to_slogic(107),
    to_slogic(109),
    to_slogic(96),
    to_slogic(92),
    to_slogic(82),
    to_slogic(96),
    to_slogic(102),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(33),
    to_slogic(33),
    to_slogic(56),
    to_slogic(102),
    to_slogic(143),
    to_slogic(170),
    to_slogic(170),
    to_slogic(170),
    to_slogic(153),
    to_slogic(133),
    to_slogic(96),
    to_slogic(44),
    to_slogic(33),
    to_slogic(89),
    to_slogic(126),
    to_slogic(152),
    to_slogic(162),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(173),
    to_slogic(156),
    to_slogic(144),
    to_slogic(117),
    to_slogic(156),
    to_slogic(91),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(50),
    to_slogic(89),
    to_slogic(120),
    to_slogic(50),
    to_slogic(56),
    to_slogic(75),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(42),
    to_slogic(83),
    to_slogic(83),
    to_slogic(83),
    to_slogic(58),
    to_slogic(65),
    to_slogic(83),
    to_slogic(89),
    to_slogic(97),
    to_slogic(115),
    to_slogic(115),
    to_slogic(76),
    to_slogic(89),
    to_slogic(91),
    to_slogic(115),
    to_slogic(136),
    to_slogic(140),
    to_slogic(138),
    to_slogic(143),
    to_slogic(75),
    to_slogic(71),
    to_slogic(42),
    to_slogic(81),
    to_slogic(153),
    to_slogic(196),
    to_slogic(102),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(75),
    to_slogic(56),
    to_slogic(75),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(97),
    to_slogic(44),
    to_slogic(44),
    to_slogic(82),
    to_slogic(109),
    to_slogic(115),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(134),
    to_slogic(134),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(149),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(177),
    to_slogic(183),
    to_slogic(183),
    to_slogic(183),
    to_slogic(187),
    to_slogic(191),
    to_slogic(198),
    to_slogic(193),
    to_slogic(207),
    to_slogic(200),
    to_slogic(211),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(220),
    to_slogic(214),
    to_slogic(220),
    to_slogic(133),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(44),
    to_slogic(36),
    to_slogic(70),
    to_slogic(143),
    to_slogic(150),
    to_slogic(137),
    to_slogic(150),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(125),
    to_slogic(124),
    to_slogic(125),
    to_slogic(118),
    to_slogic(130),
    to_slogic(157),
    to_slogic(172),
    to_slogic(183),
    to_slogic(191),
    to_slogic(205),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(203),
    to_slogic(191),
    to_slogic(136),
    to_slogic(89),
    to_slogic(82),
    to_slogic(92),
    to_slogic(96),
    to_slogic(82),
    to_slogic(96),
    to_slogic(102),
    to_slogic(101),
    to_slogic(116),
    to_slogic(116),
    to_slogic(109),
    to_slogic(94),
    to_slogic(82),
    to_slogic(92),
    to_slogic(94),
    to_slogic(101),
    to_slogic(110),
    to_slogic(96),
    to_slogic(101),
    to_slogic(33),
    to_slogic(42),
    to_slogic(49),
    to_slogic(95),
    to_slogic(149),
    to_slogic(162),
    to_slogic(170),
    to_slogic(170),
    to_slogic(165),
    to_slogic(149),
    to_slogic(91),
    to_slogic(33),
    to_slogic(44),
    to_slogic(89),
    to_slogic(135),
    to_slogic(151),
    to_slogic(165),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(172),
    to_slogic(156),
    to_slogic(151),
    to_slogic(118),
    to_slogic(109),
    to_slogic(133),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(102),
    to_slogic(127),
    to_slogic(42),
    to_slogic(49),
    to_slogic(81),
    to_slogic(49),
    to_slogic(36),
    to_slogic(50),
    to_slogic(42),
    to_slogic(63),
    to_slogic(81),
    to_slogic(89),
    to_slogic(71),
    to_slogic(58),
    to_slogic(71),
    to_slogic(91),
    to_slogic(91),
    to_slogic(107),
    to_slogic(102),
    to_slogic(89),
    to_slogic(84),
    to_slogic(84),
    to_slogic(102),
    to_slogic(145),
    to_slogic(153),
    to_slogic(145),
    to_slogic(153),
    to_slogic(81),
    to_slogic(42),
    to_slogic(71),
    to_slogic(65),
    to_slogic(168),
    to_slogic(197),
    to_slogic(81),
    to_slogic(40),
    to_slogic(36),
    to_slogic(40),
    to_slogic(75),
    to_slogic(49),
    to_slogic(83),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(92),
    to_slogic(109),
    to_slogic(109),
    to_slogic(97),
    to_slogic(100),
    to_slogic(56),
    to_slogic(49),
    to_slogic(82),
    to_slogic(109),
    to_slogic(121),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(135),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(172),
    to_slogic(177),
    to_slogic(177),
    to_slogic(177),
    to_slogic(187),
    to_slogic(183),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(205),
    to_slogic(200),
    to_slogic(200),
    to_slogic(207),
    to_slogic(204),
    to_slogic(214),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(220),
    to_slogic(195),
    to_slogic(69),
    to_slogic(44),
    to_slogic(33),
    to_slogic(44),
    to_slogic(33),
    to_slogic(75),
    to_slogic(152),
    to_slogic(143),
    to_slogic(137),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(119),
    to_slogic(125),
    to_slogic(118),
    to_slogic(124),
    to_slogic(157),
    to_slogic(178),
    to_slogic(191),
    to_slogic(191),
    to_slogic(197),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(207),
    to_slogic(196),
    to_slogic(169),
    to_slogic(116),
    to_slogic(94),
    to_slogic(82),
    to_slogic(100),
    to_slogic(92),
    to_slogic(96),
    to_slogic(100),
    to_slogic(101),
    to_slogic(109),
    to_slogic(107),
    to_slogic(109),
    to_slogic(96),
    to_slogic(92),
    to_slogic(94),
    to_slogic(92),
    to_slogic(101),
    to_slogic(109),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(33),
    to_slogic(40),
    to_slogic(49),
    to_slogic(89),
    to_slogic(149),
    to_slogic(162),
    to_slogic(170),
    to_slogic(176),
    to_slogic(165),
    to_slogic(143),
    to_slogic(88),
    to_slogic(33),
    to_slogic(44),
    to_slogic(89),
    to_slogic(130),
    to_slogic(152),
    to_slogic(162),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(172),
    to_slogic(165),
    to_slogic(144),
    to_slogic(133),
    to_slogic(126),
    to_slogic(119),
    to_slogic(49),
    to_slogic(56),
    to_slogic(42),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(58),
    to_slogic(130),
    to_slogic(119),
    to_slogic(49),
    to_slogic(42),
    to_slogic(68),
    to_slogic(63),
    to_slogic(40),
    to_slogic(63),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(78),
    to_slogic(76),
    to_slogic(97),
    to_slogic(102),
    to_slogic(97),
    to_slogic(84),
    to_slogic(84),
    to_slogic(78),
    to_slogic(103),
    to_slogic(138),
    to_slogic(145),
    to_slogic(120),
    to_slogic(162),
    to_slogic(107),
    to_slogic(49),
    to_slogic(50),
    to_slogic(56),
    to_slogic(168),
    to_slogic(177),
    to_slogic(68),
    to_slogic(40),
    to_slogic(40),
    to_slogic(56),
    to_slogic(82),
    to_slogic(56),
    to_slogic(88),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(70),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(56),
    to_slogic(56),
    to_slogic(83),
    to_slogic(102),
    to_slogic(118),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(134),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(144),
    to_slogic(152),
    to_slogic(149),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(187),
    to_slogic(183),
    to_slogic(183),
    to_slogic(187),
    to_slogic(191),
    to_slogic(193),
    to_slogic(198),
    to_slogic(200),
    to_slogic(207),
    to_slogic(211),
    to_slogic(204),
    to_slogic(213),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(214),
    to_slogic(125),
    to_slogic(33),
    to_slogic(33),
    to_slogic(33),
    to_slogic(36),
    to_slogic(92),
    to_slogic(152),
    to_slogic(150),
    to_slogic(137),
    to_slogic(143),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(124),
    to_slogic(125),
    to_slogic(130),
    to_slogic(144),
    to_slogic(178),
    to_slogic(191),
    to_slogic(197),
    to_slogic(197),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(203),
    to_slogic(184),
    to_slogic(144),
    to_slogic(100),
    to_slogic(92),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(94),
    to_slogic(101),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(96),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(109),
    to_slogic(101),
    to_slogic(96),
    to_slogic(101),
    to_slogic(109),
    to_slogic(33),
    to_slogic(33),
    to_slogic(49),
    to_slogic(91),
    to_slogic(127),
    to_slogic(153),
    to_slogic(170),
    to_slogic(170),
    to_slogic(165),
    to_slogic(133),
    to_slogic(96),
    to_slogic(33),
    to_slogic(44),
    to_slogic(89),
    to_slogic(121),
    to_slogic(156),
    to_slogic(165),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(172),
    to_slogic(157),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(89),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(83),
    to_slogic(138),
    to_slogic(102),
    to_slogic(40),
    to_slogic(40),
    to_slogic(56),
    to_slogic(63),
    to_slogic(40),
    to_slogic(68),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(42),
    to_slogic(56),
    to_slogic(50),
    to_slogic(81),
    to_slogic(65),
    to_slogic(97),
    to_slogic(102),
    to_slogic(107),
    to_slogic(97),
    to_slogic(78),
    to_slogic(71),
    to_slogic(107),
    to_slogic(145),
    to_slogic(120),
    to_slogic(136),
    to_slogic(153),
    to_slogic(120),
    to_slogic(81),
    to_slogic(42),
    to_slogic(56),
    to_slogic(168),
    to_slogic(127),
    to_slogic(71),
    to_slogic(42),
    to_slogic(36),
    to_slogic(56),
    to_slogic(82),
    to_slogic(56),
    to_slogic(75),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(92),
    to_slogic(100),
    to_slogic(115),
    to_slogic(124),
    to_slogic(109),
    to_slogic(56),
    to_slogic(49),
    to_slogic(92),
    to_slogic(109),
    to_slogic(121),
    to_slogic(134),
    to_slogic(124),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(130),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(162),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(177),
    to_slogic(176),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(198),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(223),
    to_slogic(176),
    to_slogic(49),
    to_slogic(33),
    to_slogic(33),
    to_slogic(33),
    to_slogic(101),
    to_slogic(144),
    to_slogic(137),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(125),
    to_slogic(130),
    to_slogic(124),
    to_slogic(118),
    to_slogic(133),
    to_slogic(173),
    to_slogic(198),
    to_slogic(213),
    to_slogic(207),
    to_slogic(205),
    to_slogic(197),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(196),
    to_slogic(175),
    to_slogic(130),
    to_slogic(89),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(107),
    to_slogic(116),
    to_slogic(96),
    to_slogic(92),
    to_slogic(83),
    to_slogic(96),
    to_slogic(109),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(109),
    to_slogic(101),
    to_slogic(33),
    to_slogic(33),
    to_slogic(36),
    to_slogic(81),
    to_slogic(133),
    to_slogic(153),
    to_slogic(170),
    to_slogic(170),
    to_slogic(170),
    to_slogic(143),
    to_slogic(88),
    to_slogic(33),
    to_slogic(44),
    to_slogic(81),
    to_slogic(126),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(184),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(161),
    to_slogic(143),
    to_slogic(144),
    to_slogic(133),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(36),
    to_slogic(50),
    to_slogic(122),
    to_slogic(127),
    to_slogic(102),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(49),
    to_slogic(50),
    to_slogic(50),
    to_slogic(63),
    to_slogic(71),
    to_slogic(84),
    to_slogic(102),
    to_slogic(120),
    to_slogic(83),
    to_slogic(65),
    to_slogic(58),
    to_slogic(97),
    to_slogic(153),
    to_slogic(136),
    to_slogic(145),
    to_slogic(127),
    to_slogic(102),
    to_slogic(138),
    to_slogic(103),
    to_slogic(107),
    to_slogic(163),
    to_slogic(102),
    to_slogic(162),
    to_slogic(68),
    to_slogic(40),
    to_slogic(64),
    to_slogic(75),
    to_slogic(56),
    to_slogic(70),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(81),
    to_slogic(115),
    to_slogic(116),
    to_slogic(126),
    to_slogic(121),
    to_slogic(109),
    to_slogic(63),
    to_slogic(56),
    to_slogic(92),
    to_slogic(109),
    to_slogic(121),
    to_slogic(130),
    to_slogic(134),
    to_slogic(134),
    to_slogic(130),
    to_slogic(139),
    to_slogic(135),
    to_slogic(134),
    to_slogic(135),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(177),
    to_slogic(177),
    to_slogic(183),
    to_slogic(183),
    to_slogic(187),
    to_slogic(191),
    to_slogic(193),
    to_slogic(198),
    to_slogic(200),
    to_slogic(204),
    to_slogic(207),
    to_slogic(211),
    to_slogic(207),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(211),
    to_slogic(83),
    to_slogic(33),
    to_slogic(33),
    to_slogic(33),
    to_slogic(117),
    to_slogic(144),
    to_slogic(137),
    to_slogic(150),
    to_slogic(150),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(130),
    to_slogic(130),
    to_slogic(143),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(132),
    to_slogic(130),
    to_slogic(130),
    to_slogic(125),
    to_slogic(125),
    to_slogic(118),
    to_slogic(143),
    to_slogic(197),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(205),
    to_slogic(207),
    to_slogic(222),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(203),
    to_slogic(184),
    to_slogic(144),
    to_slogic(109),
    to_slogic(94),
    to_slogic(89),
    to_slogic(92),
    to_slogic(92),
    to_slogic(94),
    to_slogic(102),
    to_slogic(116),
    to_slogic(107),
    to_slogic(116),
    to_slogic(109),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(109),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(91),
    to_slogic(33),
    to_slogic(33),
    to_slogic(33),
    to_slogic(68),
    to_slogic(119),
    to_slogic(153),
    to_slogic(170),
    to_slogic(170),
    to_slogic(165),
    to_slogic(149),
    to_slogic(96),
    to_slogic(33),
    to_slogic(33),
    to_slogic(81),
    to_slogic(130),
    to_slogic(151),
    to_slogic(165),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(176),
    to_slogic(172),
    to_slogic(156),
    to_slogic(143),
    to_slogic(135),
    to_slogic(119),
    to_slogic(49),
    to_slogic(50),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(42),
    to_slogic(40),
    to_slogic(44),
    to_slogic(97),
    to_slogic(115),
    to_slogic(114),
    to_slogic(81),
    to_slogic(42),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(68),
    to_slogic(56),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(63),
    to_slogic(50),
    to_slogic(50),
    to_slogic(71),
    to_slogic(58),
    to_slogic(71),
    to_slogic(130),
    to_slogic(97),
    to_slogic(58),
    to_slogic(78),
    to_slogic(109),
    to_slogic(140),
    to_slogic(140),
    to_slogic(153),
    to_slogic(145),
    to_slogic(89),
    to_slogic(127),
    to_slogic(81),
    to_slogic(153),
    to_slogic(163),
    to_slogic(127),
    to_slogic(153),
    to_slogic(63),
    to_slogic(40),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(70),
    to_slogic(109),
    to_slogic(116),
    to_slogic(124),
    to_slogic(124),
    to_slogic(121),
    to_slogic(109),
    to_slogic(56),
    to_slogic(70),
    to_slogic(92),
    to_slogic(109),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(135),
    to_slogic(130),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(146),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(172),
    to_slogic(172),
    to_slogic(177),
    to_slogic(176),
    to_slogic(183),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(213),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(223),
    to_slogic(133),
    to_slogic(33),
    to_slogic(33),
    to_slogic(33),
    to_slogic(118),
    to_slogic(144),
    to_slogic(137),
    to_slogic(156),
    to_slogic(143),
    to_slogic(150),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(130),
    to_slogic(132),
    to_slogic(130),
    to_slogic(130),
    to_slogic(119),
    to_slogic(125),
    to_slogic(124),
    to_slogic(118),
    to_slogic(158),
    to_slogic(197),
    to_slogic(213),
    to_slogic(223),
    to_slogic(213),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(203),
    to_slogic(169),
    to_slogic(130),
    to_slogic(100),
    to_slogic(97),
    to_slogic(94),
    to_slogic(89),
    to_slogic(89),
    to_slogic(94),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(109),
    to_slogic(96),
    to_slogic(96),
    to_slogic(82),
    to_slogic(96),
    to_slogic(109),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(109),
    to_slogic(83),
    to_slogic(33),
    to_slogic(33),
    to_slogic(40),
    to_slogic(68),
    to_slogic(119),
    to_slogic(153),
    to_slogic(170),
    to_slogic(176),
    to_slogic(170),
    to_slogic(149),
    to_slogic(102),
    to_slogic(49),
    to_slogic(33),
    to_slogic(76),
    to_slogic(126),
    to_slogic(151),
    to_slogic(165),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(172),
    to_slogic(165),
    to_slogic(144),
    to_slogic(134),
    to_slogic(109),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(44),
    to_slogic(95),
    to_slogic(102),
    to_slogic(63),
    to_slogic(102),
    to_slogic(71),
    to_slogic(56),
    to_slogic(42),
    to_slogic(49),
    to_slogic(56),
    to_slogic(71),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(50),
    to_slogic(63),
    to_slogic(50),
    to_slogic(49),
    to_slogic(71),
    to_slogic(58),
    to_slogic(84),
    to_slogic(115),
    to_slogic(109),
    to_slogic(97),
    to_slogic(97),
    to_slogic(115),
    to_slogic(138),
    to_slogic(138),
    to_slogic(127),
    to_slogic(120),
    to_slogic(136),
    to_slogic(140),
    to_slogic(143),
    to_slogic(168),
    to_slogic(114),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(64),
    to_slogic(89),
    to_slogic(116),
    to_slogic(121),
    to_slogic(124),
    to_slogic(124),
    to_slogic(121),
    to_slogic(97),
    to_slogic(44),
    to_slogic(75),
    to_slogic(96),
    to_slogic(115),
    to_slogic(121),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(162),
    to_slogic(173),
    to_slogic(172),
    to_slogic(177),
    to_slogic(177),
    to_slogic(183),
    to_slogic(182),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(207),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(182),
    to_slogic(33),
    to_slogic(33),
    to_slogic(44),
    to_slogic(130),
    to_slogic(137),
    to_slogic(143),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(130),
    to_slogic(143),
    to_slogic(132),
    to_slogic(130),
    to_slogic(132),
    to_slogic(130),
    to_slogic(125),
    to_slogic(124),
    to_slogic(118),
    to_slogic(124),
    to_slogic(158),
    to_slogic(207),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(205),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(203),
    to_slogic(184),
    to_slogic(156),
    to_slogic(118),
    to_slogic(109),
    to_slogic(100),
    to_slogic(100),
    to_slogic(89),
    to_slogic(94),
    to_slogic(100),
    to_slogic(102),
    to_slogic(116),
    to_slogic(109),
    to_slogic(102),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(109),
    to_slogic(101),
    to_slogic(110),
    to_slogic(101),
    to_slogic(91),
    to_slogic(101),
    to_slogic(83),
    to_slogic(83),
    to_slogic(33),
    to_slogic(33),
    to_slogic(36),
    to_slogic(68),
    to_slogic(119),
    to_slogic(153),
    to_slogic(170),
    to_slogic(170),
    to_slogic(170),
    to_slogic(143),
    to_slogic(102),
    to_slogic(49),
    to_slogic(44),
    to_slogic(81),
    to_slogic(126),
    to_slogic(152),
    to_slogic(165),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(165),
    to_slogic(157),
    to_slogic(152),
    to_slogic(133),
    to_slogic(113),
    to_slogic(69),
    to_slogic(63),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(71),
    to_slogic(68),
    to_slogic(50),
    to_slogic(63),
    to_slogic(107),
    to_slogic(81),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(68),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(63),
    to_slogic(50),
    to_slogic(42),
    to_slogic(89),
    to_slogic(56),
    to_slogic(50),
    to_slogic(71),
    to_slogic(89),
    to_slogic(122),
    to_slogic(130),
    to_slogic(122),
    to_slogic(130),
    to_slogic(143),
    to_slogic(102),
    to_slogic(81),
    to_slogic(120),
    to_slogic(130),
    to_slogic(163),
    to_slogic(153),
    to_slogic(138),
    to_slogic(89),
    to_slogic(63),
    to_slogic(91),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(76),
    to_slogic(89),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(124),
    to_slogic(117),
    to_slogic(97),
    to_slogic(44),
    to_slogic(81),
    to_slogic(92),
    to_slogic(115),
    to_slogic(124),
    to_slogic(130),
    to_slogic(134),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(144),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(176),
    to_slogic(177),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(214),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(220),
    to_slogic(211),
    to_slogic(64),
    to_slogic(33),
    to_slogic(40),
    to_slogic(137),
    to_slogic(136),
    to_slogic(143),
    to_slogic(143),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(130),
    to_slogic(132),
    to_slogic(132),
    to_slogic(119),
    to_slogic(130),
    to_slogic(124),
    to_slogic(118),
    to_slogic(133),
    to_slogic(178),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(205),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(203),
    to_slogic(175),
    to_slogic(136),
    to_slogic(121),
    to_slogic(109),
    to_slogic(102),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(107),
    to_slogic(102),
    to_slogic(96),
    to_slogic(92),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(96),
    to_slogic(83),
    to_slogic(83),
    to_slogic(33),
    to_slogic(33),
    to_slogic(33),
    to_slogic(63),
    to_slogic(113),
    to_slogic(153),
    to_slogic(162),
    to_slogic(170),
    to_slogic(170),
    to_slogic(149),
    to_slogic(119),
    to_slogic(62),
    to_slogic(33),
    to_slogic(75),
    to_slogic(121),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(157),
    to_slogic(144),
    to_slogic(133),
    to_slogic(133),
    to_slogic(71),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(89),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(81),
    to_slogic(89),
    to_slogic(63),
    to_slogic(49),
    to_slogic(42),
    to_slogic(68),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(50),
    to_slogic(68),
    to_slogic(50),
    to_slogic(56),
    to_slogic(89),
    to_slogic(65),
    to_slogic(49),
    to_slogic(42),
    to_slogic(58),
    to_slogic(107),
    to_slogic(140),
    to_slogic(130),
    to_slogic(120),
    to_slogic(138),
    to_slogic(115),
    to_slogic(102),
    to_slogic(68),
    to_slogic(81),
    to_slogic(113),
    to_slogic(114),
    to_slogic(143),
    to_slogic(133),
    to_slogic(127),
    to_slogic(113),
    to_slogic(102),
    to_slogic(95),
    to_slogic(63),
    to_slogic(75),
    to_slogic(64),
    to_slogic(83),
    to_slogic(82),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(76),
    to_slogic(75),
    to_slogic(100),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(124),
    to_slogic(124),
    to_slogic(89),
    to_slogic(56),
    to_slogic(82),
    to_slogic(96),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(149),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(173),
    to_slogic(165),
    to_slogic(177),
    to_slogic(183),
    to_slogic(182),
    to_slogic(191),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(213),
    to_slogic(109),
    to_slogic(33),
    to_slogic(62),
    to_slogic(130),
    to_slogic(137),
    to_slogic(143),
    to_slogic(150),
    to_slogic(156),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(130),
    to_slogic(143),
    to_slogic(132),
    to_slogic(130),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(119),
    to_slogic(124),
    to_slogic(124),
    to_slogic(136),
    to_slogic(183),
    to_slogic(207),
    to_slogic(213),
    to_slogic(207),
    to_slogic(205),
    to_slogic(205),
    to_slogic(207),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(203),
    to_slogic(184),
    to_slogic(144),
    to_slogic(130),
    to_slogic(116),
    to_slogic(116),
    to_slogic(100),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(102),
    to_slogic(102),
    to_slogic(116),
    to_slogic(109),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(109),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(101),
    to_slogic(83),
    to_slogic(87),
    to_slogic(83),
    to_slogic(33),
    to_slogic(33),
    to_slogic(36),
    to_slogic(63),
    to_slogic(114),
    to_slogic(153),
    to_slogic(170),
    to_slogic(170),
    to_slogic(170),
    to_slogic(153),
    to_slogic(118),
    to_slogic(49),
    to_slogic(44),
    to_slogic(76),
    to_slogic(121),
    to_slogic(151),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(165),
    to_slogic(156),
    to_slogic(144),
    to_slogic(149),
    to_slogic(121),
    to_slogic(75),
    to_slogic(56),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(89),
    to_slogic(68),
    to_slogic(63),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(68),
    to_slogic(44),
    to_slogic(71),
    to_slogic(95),
    to_slogic(49),
    to_slogic(50),
    to_slogic(44),
    to_slogic(58),
    to_slogic(97),
    to_slogic(138),
    to_slogic(115),
    to_slogic(140),
    to_slogic(115),
    to_slogic(127),
    to_slogic(95),
    to_slogic(63),
    to_slogic(33),
    to_slogic(68),
    to_slogic(68),
    to_slogic(49),
    to_slogic(64),
    to_slogic(82),
    to_slogic(68),
    to_slogic(102),
    to_slogic(114),
    to_slogic(113),
    to_slogic(143),
    to_slogic(113),
    to_slogic(91),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(70),
    to_slogic(92),
    to_slogic(109),
    to_slogic(117),
    to_slogic(121),
    to_slogic(130),
    to_slogic(126),
    to_slogic(121),
    to_slogic(82),
    to_slogic(56),
    to_slogic(82),
    to_slogic(109),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(130),
    to_slogic(139),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(162),
    to_slogic(177),
    to_slogic(177),
    to_slogic(187),
    to_slogic(182),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(200),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(223),
    to_slogic(162),
    to_slogic(36),
    to_slogic(75),
    to_slogic(130),
    to_slogic(144),
    to_slogic(143),
    to_slogic(150),
    to_slogic(150),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(119),
    to_slogic(130),
    to_slogic(124),
    to_slogic(124),
    to_slogic(137),
    to_slogic(183),
    to_slogic(207),
    to_slogic(213),
    to_slogic(213),
    to_slogic(205),
    to_slogic(205),
    to_slogic(207),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(203),
    to_slogic(175),
    to_slogic(136),
    to_slogic(121),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(94),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(94),
    to_slogic(94),
    to_slogic(89),
    to_slogic(92),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(91),
    to_slogic(96),
    to_slogic(83),
    to_slogic(96),
    to_slogic(91),
    to_slogic(36),
    to_slogic(33),
    to_slogic(33),
    to_slogic(56),
    to_slogic(95),
    to_slogic(153),
    to_slogic(165),
    to_slogic(170),
    to_slogic(176),
    to_slogic(156),
    to_slogic(119),
    to_slogic(49),
    to_slogic(44),
    to_slogic(75),
    to_slogic(121),
    to_slogic(151),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(172),
    to_slogic(165),
    to_slogic(144),
    to_slogic(151),
    to_slogic(101),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(71),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(68),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(42),
    to_slogic(63),
    to_slogic(42),
    to_slogic(81),
    to_slogic(95),
    to_slogic(42),
    to_slogic(71),
    to_slogic(58),
    to_slogic(71),
    to_slogic(97),
    to_slogic(115),
    to_slogic(102),
    to_slogic(130),
    to_slogic(107),
    to_slogic(115),
    to_slogic(120),
    to_slogic(115),
    to_slogic(49),
    to_slogic(56),
    to_slogic(81),
    to_slogic(33),
    to_slogic(64),
    to_slogic(40),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(64),
    to_slogic(88),
    to_slogic(64),
    to_slogic(102),
    to_slogic(96),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(89),
    to_slogic(89),
    to_slogic(115),
    to_slogic(121),
    to_slogic(126),
    to_slogic(130),
    to_slogic(128),
    to_slogic(121),
    to_slogic(70),
    to_slogic(63),
    to_slogic(92),
    to_slogic(102),
    to_slogic(124),
    to_slogic(134),
    to_slogic(130),
    to_slogic(134),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(151),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(173),
    to_slogic(165),
    to_slogic(172),
    to_slogic(177),
    to_slogic(177),
    to_slogic(183),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(214),
    to_slogic(213),
    to_slogic(193),
    to_slogic(49),
    to_slogic(82),
    to_slogic(130),
    to_slogic(137),
    to_slogic(143),
    to_slogic(150),
    to_slogic(150),
    to_slogic(156),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(130),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(130),
    to_slogic(119),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(136),
    to_slogic(183),
    to_slogic(205),
    to_slogic(213),
    to_slogic(205),
    to_slogic(205),
    to_slogic(205),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(203),
    to_slogic(196),
    to_slogic(161),
    to_slogic(130),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(102),
    to_slogic(100),
    to_slogic(92),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(100),
    to_slogic(92),
    to_slogic(82),
    to_slogic(89),
    to_slogic(96),
    to_slogic(101),
    to_slogic(110),
    to_slogic(101),
    to_slogic(96),
    to_slogic(96),
    to_slogic(96),
    to_slogic(87),
    to_slogic(91),
    to_slogic(91),
    to_slogic(33),
    to_slogic(33),
    to_slogic(40),
    to_slogic(49),
    to_slogic(102),
    to_slogic(143),
    to_slogic(162),
    to_slogic(176),
    to_slogic(170),
    to_slogic(153),
    to_slogic(119),
    to_slogic(64),
    to_slogic(49),
    to_slogic(75),
    to_slogic(116),
    to_slogic(144),
    to_slogic(165),
    to_slogic(172),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(172),
    to_slogic(165),
    to_slogic(144),
    to_slogic(155),
    to_slogic(110),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(42),
    to_slogic(40),
    to_slogic(42),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(68),
    to_slogic(49),
    to_slogic(50),
    to_slogic(50),
    to_slogic(68),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(68),
    to_slogic(63),
    to_slogic(40),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(44),
    to_slogic(83),
    to_slogic(71),
    to_slogic(76),
    to_slogic(50),
    to_slogic(91),
    to_slogic(83),
    to_slogic(97),
    to_slogic(102),
    to_slogic(120),
    to_slogic(107),
    to_slogic(115),
    to_slogic(107),
    to_slogic(122),
    to_slogic(138),
    to_slogic(89),
    to_slogic(56),
    to_slogic(95),
    to_slogic(40),
    to_slogic(56),
    to_slogic(40),
    to_slogic(56),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(88),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(62),
    to_slogic(75),
    to_slogic(89),
    to_slogic(100),
    to_slogic(116),
    to_slogic(124),
    to_slogic(124),
    to_slogic(128),
    to_slogic(126),
    to_slogic(109),
    to_slogic(70),
    to_slogic(70),
    to_slogic(96),
    to_slogic(117),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(182),
    to_slogic(183),
    to_slogic(193),
    to_slogic(193),
    to_slogic(189),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(204),
    to_slogic(87),
    to_slogic(92),
    to_slogic(130),
    to_slogic(143),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(133),
    to_slogic(132),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(132),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(137),
    to_slogic(165),
    to_slogic(191),
    to_slogic(205),
    to_slogic(203),
    to_slogic(196),
    to_slogic(205),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(213),
    to_slogic(191),
    to_slogic(144),
    to_slogic(121),
    to_slogic(116),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(94),
    to_slogic(94),
    to_slogic(99),
    to_slogic(96),
    to_slogic(100),
    to_slogic(92),
    to_slogic(75),
    to_slogic(92),
    to_slogic(96),
    to_slogic(109),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(91),
    to_slogic(96),
    to_slogic(91),
    to_slogic(91),
    to_slogic(96),
    to_slogic(96),
    to_slogic(33),
    to_slogic(40),
    to_slogic(33),
    to_slogic(42),
    to_slogic(96),
    to_slogic(149),
    to_slogic(153),
    to_slogic(170),
    to_slogic(170),
    to_slogic(165),
    to_slogic(119),
    to_slogic(64),
    to_slogic(49),
    to_slogic(76),
    to_slogic(116),
    to_slogic(151),
    to_slogic(157),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(172),
    to_slogic(157),
    to_slogic(144),
    to_slogic(157),
    to_slogic(127),
    to_slogic(69),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(81),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(50),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(50),
    to_slogic(63),
    to_slogic(89),
    to_slogic(63),
    to_slogic(95),
    to_slogic(71),
    to_slogic(63),
    to_slogic(109),
    to_slogic(91),
    to_slogic(97),
    to_slogic(115),
    to_slogic(130),
    to_slogic(115),
    to_slogic(71),
    to_slogic(89),
    to_slogic(120),
    to_slogic(130),
    to_slogic(75),
    to_slogic(89),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(62),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(92),
    to_slogic(109),
    to_slogic(115),
    to_slogic(124),
    to_slogic(126),
    to_slogic(130),
    to_slogic(126),
    to_slogic(100),
    to_slogic(63),
    to_slogic(82),
    to_slogic(96),
    to_slogic(116),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(155),
    to_slogic(161),
    to_slogic(162),
    to_slogic(162),
    to_slogic(173),
    to_slogic(165),
    to_slogic(166),
    to_slogic(183),
    to_slogic(183),
    to_slogic(183),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(214),
    to_slogic(213),
    to_slogic(133),
    to_slogic(92),
    to_slogic(130),
    to_slogic(144),
    to_slogic(143),
    to_slogic(150),
    to_slogic(150),
    to_slogic(149),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(133),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(132),
    to_slogic(130),
    to_slogic(132),
    to_slogic(137),
    to_slogic(124),
    to_slogic(137),
    to_slogic(136),
    to_slogic(144),
    to_slogic(169),
    to_slogic(184),
    to_slogic(191),
    to_slogic(191),
    to_slogic(205),
    to_slogic(213),
    to_slogic(213),
    to_slogic(213),
    to_slogic(203),
    to_slogic(175),
    to_slogic(143),
    to_slogic(121),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(89),
    to_slogic(92),
    to_slogic(94),
    to_slogic(109),
    to_slogic(82),
    to_slogic(76),
    to_slogic(81),
    to_slogic(96),
    to_slogic(101),
    to_slogic(109),
    to_slogic(96),
    to_slogic(101),
    to_slogic(83),
    to_slogic(96),
    to_slogic(96),
    to_slogic(91),
    to_slogic(101),
    to_slogic(91),
    to_slogic(91),
    to_slogic(40),
    to_slogic(40),
    to_slogic(36),
    to_slogic(49),
    to_slogic(81),
    to_slogic(133),
    to_slogic(162),
    to_slogic(170),
    to_slogic(170),
    to_slogic(153),
    to_slogic(119),
    to_slogic(88),
    to_slogic(49),
    to_slogic(75),
    to_slogic(121),
    to_slogic(143),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(165),
    to_slogic(165),
    to_slogic(144),
    to_slogic(155),
    to_slogic(133),
    to_slogic(69),
    to_slogic(81),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(50),
    to_slogic(63),
    to_slogic(81),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(68),
    to_slogic(63),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(50),
    to_slogic(81),
    to_slogic(49),
    to_slogic(50),
    to_slogic(49),
    to_slogic(71),
    to_slogic(71),
    to_slogic(63),
    to_slogic(65),
    to_slogic(71),
    to_slogic(95),
    to_slogic(44),
    to_slogic(71),
    to_slogic(145),
    to_slogic(130),
    to_slogic(132),
    to_slogic(120),
    to_slogic(102),
    to_slogic(89),
    to_slogic(65),
    to_slogic(102),
    to_slogic(122),
    to_slogic(122),
    to_slogic(107),
    to_slogic(115),
    to_slogic(81),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(75),
    to_slogic(89),
    to_slogic(89),
    to_slogic(109),
    to_slogic(116),
    to_slogic(124),
    to_slogic(124),
    to_slogic(126),
    to_slogic(121),
    to_slogic(82),
    to_slogic(56),
    to_slogic(83),
    to_slogic(109),
    to_slogic(117),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(139),
    to_slogic(139),
    to_slogic(134),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(130),
    to_slogic(139),
    to_slogic(135),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(146),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(162),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(177),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(213),
    to_slogic(176),
    to_slogic(116),
    to_slogic(136),
    to_slogic(143),
    to_slogic(124),
    to_slogic(130),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(143),
    to_slogic(149),
    to_slogic(150),
    to_slogic(150),
    to_slogic(144),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(132),
    to_slogic(130),
    to_slogic(130),
    to_slogic(144),
    to_slogic(137),
    to_slogic(136),
    to_slogic(136),
    to_slogic(144),
    to_slogic(161),
    to_slogic(161),
    to_slogic(184),
    to_slogic(207),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(203),
    to_slogic(175),
    to_slogic(130),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(100),
    to_slogic(99),
    to_slogic(92),
    to_slogic(94),
    to_slogic(102),
    to_slogic(92),
    to_slogic(89),
    to_slogic(75),
    to_slogic(82),
    to_slogic(109),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(96),
    to_slogic(83),
    to_slogic(96),
    to_slogic(91),
    to_slogic(96),
    to_slogic(96),
    to_slogic(101),
    to_slogic(83),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(42),
    to_slogic(68),
    to_slogic(133),
    to_slogic(153),
    to_slogic(170),
    to_slogic(170),
    to_slogic(166),
    to_slogic(133),
    to_slogic(91),
    to_slogic(56),
    to_slogic(76),
    to_slogic(116),
    to_slogic(144),
    to_slogic(165),
    to_slogic(172),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(157),
    to_slogic(144),
    to_slogic(152),
    to_slogic(141),
    to_slogic(75),
    to_slogic(81),
    to_slogic(56),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(68),
    to_slogic(81),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(50),
    to_slogic(63),
    to_slogic(63),
    to_slogic(68),
    to_slogic(63),
    to_slogic(49),
    to_slogic(63),
    to_slogic(64),
    to_slogic(56),
    to_slogic(42),
    to_slogic(81),
    to_slogic(83),
    to_slogic(42),
    to_slogic(49),
    to_slogic(63),
    to_slogic(102),
    to_slogic(71),
    to_slogic(50),
    to_slogic(68),
    to_slogic(81),
    to_slogic(102),
    to_slogic(120),
    to_slogic(115),
    to_slogic(71),
    to_slogic(50),
    to_slogic(76),
    to_slogic(117),
    to_slogic(145),
    to_slogic(145),
    to_slogic(162),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(62),
    to_slogic(75),
    to_slogic(89),
    to_slogic(109),
    to_slogic(115),
    to_slogic(121),
    to_slogic(126),
    to_slogic(124),
    to_slogic(126),
    to_slogic(109),
    to_slogic(70),
    to_slogic(64),
    to_slogic(92),
    to_slogic(117),
    to_slogic(130),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(130),
    to_slogic(139),
    to_slogic(130),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(155),
    to_slogic(165),
    to_slogic(178),
    to_slogic(166),
    to_slogic(183),
    to_slogic(183),
    to_slogic(182),
    to_slogic(193),
    to_slogic(193),
    to_slogic(198),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(200),
    to_slogic(133),
    to_slogic(144),
    to_slogic(136),
    to_slogic(107),
    to_slogic(118),
    to_slogic(118),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(130),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(143),
    to_slogic(136),
    to_slogic(130),
    to_slogic(144),
    to_slogic(184),
    to_slogic(205),
    to_slogic(222),
    to_slogic(222),
    to_slogic(203),
    to_slogic(196),
    to_slogic(161),
    to_slogic(130),
    to_slogic(116),
    to_slogic(109),
    to_slogic(100),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(96),
    to_slogic(100),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(96),
    to_slogic(109),
    to_slogic(101),
    to_slogic(96),
    to_slogic(96),
    to_slogic(92),
    to_slogic(87),
    to_slogic(91),
    to_slogic(96),
    to_slogic(91),
    to_slogic(96),
    to_slogic(91),
    to_slogic(75),
    to_slogic(33),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(81),
    to_slogic(133),
    to_slogic(153),
    to_slogic(170),
    to_slogic(165),
    to_slogic(153),
    to_slogic(133),
    to_slogic(88),
    to_slogic(56),
    to_slogic(75),
    to_slogic(116),
    to_slogic(143),
    to_slogic(157),
    to_slogic(172),
    to_slogic(173),
    to_slogic(176),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(172),
    to_slogic(157),
    to_slogic(144),
    to_slogic(144),
    to_slogic(141),
    to_slogic(68),
    to_slogic(87),
    to_slogic(56),
    to_slogic(42),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(42),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(89),
    to_slogic(63),
    to_slogic(42),
    to_slogic(44),
    to_slogic(76),
    to_slogic(120),
    to_slogic(84),
    to_slogic(71),
    to_slogic(49),
    to_slogic(56),
    to_slogic(50),
    to_slogic(81),
    to_slogic(138),
    to_slogic(83),
    to_slogic(50),
    to_slogic(76),
    to_slogic(81),
    to_slogic(113),
    to_slogic(162),
    to_slogic(102),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(100),
    to_slogic(109),
    to_slogic(116),
    to_slogic(121),
    to_slogic(124),
    to_slogic(121),
    to_slogic(121),
    to_slogic(99),
    to_slogic(49),
    to_slogic(75),
    to_slogic(100),
    to_slogic(121),
    to_slogic(130),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(135),
    to_slogic(134),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(146),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(177),
    to_slogic(177),
    to_slogic(183),
    to_slogic(187),
    to_slogic(193),
    to_slogic(189),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(155),
    to_slogic(143),
    to_slogic(118),
    to_slogic(94),
    to_slogic(88),
    to_slogic(102),
    to_slogic(102),
    to_slogic(107),
    to_slogic(118),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(149),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(130),
    to_slogic(143),
    to_slogic(143),
    to_slogic(144),
    to_slogic(143),
    to_slogic(144),
    to_slogic(136),
    to_slogic(136),
    to_slogic(136),
    to_slogic(157),
    to_slogic(191),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(203),
    to_slogic(184),
    to_slogic(156),
    to_slogic(121),
    to_slogic(109),
    to_slogic(109),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(92),
    to_slogic(100),
    to_slogic(92),
    to_slogic(75),
    to_slogic(75),
    to_slogic(92),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(91),
    to_slogic(83),
    to_slogic(96),
    to_slogic(96),
    to_slogic(101),
    to_slogic(91),
    to_slogic(91),
    to_slogic(82),
    to_slogic(64),
    to_slogic(40),
    to_slogic(33),
    to_slogic(33),
    to_slogic(40),
    to_slogic(68),
    to_slogic(119),
    to_slogic(153),
    to_slogic(162),
    to_slogic(176),
    to_slogic(165),
    to_slogic(133),
    to_slogic(91),
    to_slogic(62),
    to_slogic(81),
    to_slogic(109),
    to_slogic(144),
    to_slogic(158),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(165),
    to_slogic(143),
    to_slogic(128),
    to_slogic(134),
    to_slogic(75),
    to_slogic(81),
    to_slogic(63),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(81),
    to_slogic(68),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(49),
    to_slogic(81),
    to_slogic(49),
    to_slogic(56),
    to_slogic(50),
    to_slogic(71),
    to_slogic(122),
    to_slogic(127),
    to_slogic(71),
    to_slogic(71),
    to_slogic(49),
    to_slogic(42),
    to_slogic(50),
    to_slogic(102),
    to_slogic(89),
    to_slogic(50),
    to_slogic(89),
    to_slogic(115),
    to_slogic(84),
    to_slogic(119),
    to_slogic(68),
    to_slogic(40),
    to_slogic(62),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(75),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(126),
    to_slogic(126),
    to_slogic(116),
    to_slogic(81),
    to_slogic(49),
    to_slogic(82),
    to_slogic(109),
    to_slogic(134),
    to_slogic(130),
    to_slogic(139),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(146),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(162),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(183),
    to_slogic(182),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(204),
    to_slogic(200),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(220),
    to_slogic(187),
    to_slogic(118),
    to_slogic(94),
    to_slogic(75),
    to_slogic(82),
    to_slogic(89),
    to_slogic(88),
    to_slogic(88),
    to_slogic(102),
    to_slogic(107),
    to_slogic(107),
    to_slogic(109),
    to_slogic(124),
    to_slogic(125),
    to_slogic(130),
    to_slogic(130),
    to_slogic(132),
    to_slogic(143),
    to_slogic(132),
    to_slogic(143),
    to_slogic(143),
    to_slogic(143),
    to_slogic(150),
    to_slogic(158),
    to_slogic(156),
    to_slogic(136),
    to_slogic(136),
    to_slogic(136),
    to_slogic(136),
    to_slogic(158),
    to_slogic(197),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(203),
    to_slogic(175),
    to_slogic(136),
    to_slogic(116),
    to_slogic(109),
    to_slogic(92),
    to_slogic(89),
    to_slogic(81),
    to_slogic(92),
    to_slogic(100),
    to_slogic(94),
    to_slogic(75),
    to_slogic(70),
    to_slogic(82),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(96),
    to_slogic(96),
    to_slogic(96),
    to_slogic(83),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(91),
    to_slogic(83),
    to_slogic(64),
    to_slogic(62),
    to_slogic(33),
    to_slogic(33),
    to_slogic(40),
    to_slogic(40),
    to_slogic(63),
    to_slogic(114),
    to_slogic(153),
    to_slogic(177),
    to_slogic(170),
    to_slogic(170),
    to_slogic(149),
    to_slogic(102),
    to_slogic(64),
    to_slogic(70),
    to_slogic(109),
    to_slogic(143),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(178),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(172),
    to_slogic(161),
    to_slogic(151),
    to_slogic(130),
    to_slogic(120),
    to_slogic(87),
    to_slogic(81),
    to_slogic(63),
    to_slogic(42),
    to_slogic(40),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(50),
    to_slogic(71),
    to_slogic(91),
    to_slogic(84),
    to_slogic(107),
    to_slogic(130),
    to_slogic(115),
    to_slogic(50),
    to_slogic(65),
    to_slogic(63),
    to_slogic(50),
    to_slogic(63),
    to_slogic(63),
    to_slogic(50),
    to_slogic(95),
    to_slogic(89),
    to_slogic(95),
    to_slogic(102),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(33),
    to_slogic(33),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(75),
    to_slogic(97),
    to_slogic(116),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(100),
    to_slogic(44),
    to_slogic(70),
    to_slogic(92),
    to_slogic(117),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(143),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(151),
    to_slogic(165),
    to_slogic(155),
    to_slogic(165),
    to_slogic(162),
    to_slogic(173),
    to_slogic(162),
    to_slogic(177),
    to_slogic(177),
    to_slogic(183),
    to_slogic(193),
    to_slogic(182),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(204),
    to_slogic(109),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(70),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(94),
    to_slogic(102),
    to_slogic(102),
    to_slogic(102),
    to_slogic(107),
    to_slogic(118),
    to_slogic(114),
    to_slogic(119),
    to_slogic(130),
    to_slogic(132),
    to_slogic(143),
    to_slogic(150),
    to_slogic(158),
    to_slogic(158),
    to_slogic(144),
    to_slogic(144),
    to_slogic(118),
    to_slogic(136),
    to_slogic(136),
    to_slogic(184),
    to_slogic(205),
    to_slogic(213),
    to_slogic(222),
    to_slogic(203),
    to_slogic(191),
    to_slogic(161),
    to_slogic(121),
    to_slogic(109),
    to_slogic(97),
    to_slogic(89),
    to_slogic(70),
    to_slogic(82),
    to_slogic(94),
    to_slogic(100),
    to_slogic(82),
    to_slogic(70),
    to_slogic(82),
    to_slogic(92),
    to_slogic(101),
    to_slogic(96),
    to_slogic(96),
    to_slogic(96),
    to_slogic(96),
    to_slogic(87),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(91),
    to_slogic(87),
    to_slogic(82),
    to_slogic(64),
    to_slogic(56),
    to_slogic(33),
    to_slogic(33),
    to_slogic(33),
    to_slogic(40),
    to_slogic(56),
    to_slogic(119),
    to_slogic(153),
    to_slogic(176),
    to_slogic(177),
    to_slogic(170),
    to_slogic(149),
    to_slogic(102),
    to_slogic(49),
    to_slogic(70),
    to_slogic(109),
    to_slogic(135),
    to_slogic(157),
    to_slogic(173),
    to_slogic(172),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(172),
    to_slogic(165),
    to_slogic(143),
    to_slogic(133),
    to_slogic(117),
    to_slogic(87),
    to_slogic(87),
    to_slogic(68),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(63),
    to_slogic(49),
    to_slogic(68),
    to_slogic(50),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(83),
    to_slogic(50),
    to_slogic(81),
    to_slogic(109),
    to_slogic(97),
    to_slogic(122),
    to_slogic(143),
    to_slogic(107),
    to_slogic(63),
    to_slogic(71),
    to_slogic(56),
    to_slogic(75),
    to_slogic(75),
    to_slogic(71),
    to_slogic(120),
    to_slogic(68),
    to_slogic(68),
    to_slogic(88),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(33),
    to_slogic(62),
    to_slogic(62),
    to_slogic(75),
    to_slogic(89),
    to_slogic(109),
    to_slogic(116),
    to_slogic(121),
    to_slogic(121),
    to_slogic(109),
    to_slogic(121),
    to_slogic(116),
    to_slogic(62),
    to_slogic(49),
    to_slogic(75),
    to_slogic(109),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(130),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(143),
    to_slogic(144),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(155),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(166),
    to_slogic(183),
    to_slogic(182),
    to_slogic(193),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(204),
    to_slogic(200),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(120),
    to_slogic(75),
    to_slogic(82),
    to_slogic(91),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(88),
    to_slogic(88),
    to_slogic(88),
    to_slogic(102),
    to_slogic(102),
    to_slogic(118),
    to_slogic(125),
    to_slogic(143),
    to_slogic(150),
    to_slogic(158),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(183),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(203),
    to_slogic(175),
    to_slogic(136),
    to_slogic(116),
    to_slogic(94),
    to_slogic(81),
    to_slogic(75),
    to_slogic(75),
    to_slogic(92),
    to_slogic(92),
    to_slogic(82),
    to_slogic(81),
    to_slogic(75),
    to_slogic(92),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(91),
    to_slogic(96),
    to_slogic(96),
    to_slogic(91),
    to_slogic(96),
    to_slogic(109),
    to_slogic(96),
    to_slogic(91),
    to_slogic(88),
    to_slogic(75),
    to_slogic(49),
    to_slogic(56),
    to_slogic(33),
    to_slogic(40),
    to_slogic(33),
    to_slogic(33),
    to_slogic(49),
    to_slogic(119),
    to_slogic(153),
    to_slogic(177),
    to_slogic(176),
    to_slogic(176),
    to_slogic(153),
    to_slogic(119),
    to_slogic(64),
    to_slogic(70),
    to_slogic(109),
    to_slogic(143),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(121),
    to_slogic(101),
    to_slogic(96),
    to_slogic(89),
    to_slogic(63),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(68),
    to_slogic(49),
    to_slogic(50),
    to_slogic(68),
    to_slogic(56),
    to_slogic(50),
    to_slogic(56),
    to_slogic(68),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(40),
    to_slogic(49),
    to_slogic(89),
    to_slogic(84),
    to_slogic(115),
    to_slogic(120),
    to_slogic(145),
    to_slogic(120),
    to_slogic(65),
    to_slogic(83),
    to_slogic(91),
    to_slogic(122),
    to_slogic(81),
    to_slogic(75),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(70),
    to_slogic(75),
    to_slogic(100),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(116),
    to_slogic(121),
    to_slogic(116),
    to_slogic(89),
    to_slogic(44),
    to_slogic(56),
    to_slogic(96),
    to_slogic(116),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(139),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(135),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(135),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(157),
    to_slogic(155),
    to_slogic(165),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(177),
    to_slogic(187),
    to_slogic(182),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(223),
    to_slogic(149),
    to_slogic(82),
    to_slogic(89),
    to_slogic(96),
    to_slogic(94),
    to_slogic(88),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(75),
    to_slogic(70),
    to_slogic(70),
    to_slogic(64),
    to_slogic(75),
    to_slogic(64),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(88),
    to_slogic(102),
    to_slogic(124),
    to_slogic(136),
    to_slogic(144),
    to_slogic(158),
    to_slogic(158),
    to_slogic(169),
    to_slogic(144),
    to_slogic(158),
    to_slogic(197),
    to_slogic(213),
    to_slogic(222),
    to_slogic(213),
    to_slogic(196),
    to_slogic(161),
    to_slogic(121),
    to_slogic(97),
    to_slogic(75),
    to_slogic(62),
    to_slogic(62),
    to_slogic(81),
    to_slogic(89),
    to_slogic(81),
    to_slogic(89),
    to_slogic(75),
    to_slogic(82),
    to_slogic(101),
    to_slogic(107),
    to_slogic(92),
    to_slogic(96),
    to_slogic(96),
    to_slogic(91),
    to_slogic(83),
    to_slogic(96),
    to_slogic(101),
    to_slogic(102),
    to_slogic(91),
    to_slogic(91),
    to_slogic(83),
    to_slogic(64),
    to_slogic(62),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(33),
    to_slogic(40),
    to_slogic(56),
    to_slogic(114),
    to_slogic(153),
    to_slogic(170),
    to_slogic(177),
    to_slogic(176),
    to_slogic(153),
    to_slogic(132),
    to_slogic(64),
    to_slogic(70),
    to_slogic(109),
    to_slogic(130),
    to_slogic(157),
    to_slogic(165),
    to_slogic(172),
    to_slogic(176),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(165),
    to_slogic(151),
    to_slogic(92),
    to_slogic(109),
    to_slogic(96),
    to_slogic(83),
    to_slogic(63),
    to_slogic(42),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(42),
    to_slogic(63),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(68),
    to_slogic(50),
    to_slogic(49),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(49),
    to_slogic(91),
    to_slogic(107),
    to_slogic(122),
    to_slogic(138),
    to_slogic(130),
    to_slogic(117),
    to_slogic(113),
    to_slogic(91),
    to_slogic(89),
    to_slogic(102),
    to_slogic(71),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(49),
    to_slogic(33),
    to_slogic(44),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(89),
    to_slogic(100),
    to_slogic(121),
    to_slogic(109),
    to_slogic(116),
    to_slogic(121),
    to_slogic(121),
    to_slogic(97),
    to_slogic(44),
    to_slogic(44),
    to_slogic(75),
    to_slogic(109),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(143),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(155),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(165),
    to_slogic(178),
    to_slogic(177),
    to_slogic(183),
    to_slogic(182),
    to_slogic(187),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(200),
    to_slogic(211),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(185),
    to_slogic(82),
    to_slogic(82),
    to_slogic(94),
    to_slogic(101),
    to_slogic(94),
    to_slogic(94),
    to_slogic(92),
    to_slogic(92),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(64),
    to_slogic(56),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(88),
    to_slogic(101),
    to_slogic(144),
    to_slogic(183),
    to_slogic(191),
    to_slogic(184),
    to_slogic(161),
    to_slogic(176),
    to_slogic(203),
    to_slogic(213),
    to_slogic(213),
    to_slogic(203),
    to_slogic(175),
    to_slogic(136),
    to_slogic(109),
    to_slogic(81),
    to_slogic(63),
    to_slogic(56),
    to_slogic(76),
    to_slogic(81),
    to_slogic(82),
    to_slogic(75),
    to_slogic(82),
    to_slogic(92),
    to_slogic(101),
    to_slogic(110),
    to_slogic(101),
    to_slogic(96),
    to_slogic(83),
    to_slogic(92),
    to_slogic(83),
    to_slogic(96),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(91),
    to_slogic(75),
    to_slogic(64),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(63),
    to_slogic(114),
    to_slogic(153),
    to_slogic(176),
    to_slogic(177),
    to_slogic(177),
    to_slogic(170),
    to_slogic(119),
    to_slogic(75),
    to_slogic(75),
    to_slogic(109),
    to_slogic(144),
    to_slogic(157),
    to_slogic(162),
    to_slogic(172),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(173),
    to_slogic(165),
    to_slogic(151),
    to_slogic(92),
    to_slogic(120),
    to_slogic(89),
    to_slogic(69),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(68),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(50),
    to_slogic(42),
    to_slogic(50),
    to_slogic(89),
    to_slogic(107),
    to_slogic(155),
    to_slogic(130),
    to_slogic(122),
    to_slogic(120),
    to_slogic(89),
    to_slogic(91),
    to_slogic(95),
    to_slogic(83),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(33),
    to_slogic(40),
    to_slogic(33),
    to_slogic(62),
    to_slogic(70),
    to_slogic(89),
    to_slogic(94),
    to_slogic(109),
    to_slogic(121),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(109),
    to_slogic(62),
    to_slogic(44),
    to_slogic(56),
    to_slogic(96),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(135),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(155),
    to_slogic(165),
    to_slogic(162),
    to_slogic(173),
    to_slogic(172),
    to_slogic(177),
    to_slogic(183),
    to_slogic(182),
    to_slogic(187),
    to_slogic(189),
    to_slogic(200),
    to_slogic(193),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(205),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(214),
    to_slogic(213),
    to_slogic(204),
    to_slogic(110),
    to_slogic(88),
    to_slogic(94),
    to_slogic(101),
    to_slogic(101),
    to_slogic(102),
    to_slogic(101),
    to_slogic(94),
    to_slogic(94),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(118),
    to_slogic(176),
    to_slogic(197),
    to_slogic(203),
    to_slogic(175),
    to_slogic(161),
    to_slogic(184),
    to_slogic(203),
    to_slogic(213),
    to_slogic(213),
    to_slogic(203),
    to_slogic(169),
    to_slogic(121),
    to_slogic(75),
    to_slogic(62),
    to_slogic(62),
    to_slogic(63),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(70),
    to_slogic(82),
    to_slogic(96),
    to_slogic(101),
    to_slogic(107),
    to_slogic(96),
    to_slogic(83),
    to_slogic(92),
    to_slogic(83),
    to_slogic(83),
    to_slogic(96),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(91),
    to_slogic(82),
    to_slogic(64),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(83),
    to_slogic(102),
    to_slogic(149),
    to_slogic(177),
    to_slogic(189),
    to_slogic(176),
    to_slogic(170),
    to_slogic(133),
    to_slogic(82),
    to_slogic(75),
    to_slogic(109),
    to_slogic(130),
    to_slogic(157),
    to_slogic(165),
    to_slogic(173),
    to_slogic(176),
    to_slogic(172),
    to_slogic(178),
    to_slogic(176),
    to_slogic(183),
    to_slogic(172),
    to_slogic(165),
    to_slogic(144),
    to_slogic(102),
    to_slogic(121),
    to_slogic(101),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(50),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(42),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(71),
    to_slogic(122),
    to_slogic(140),
    to_slogic(138),
    to_slogic(122),
    to_slogic(91),
    to_slogic(107),
    to_slogic(102),
    to_slogic(113),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(75),
    to_slogic(75),
    to_slogic(89),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(109),
    to_slogic(76),
    to_slogic(44),
    to_slogic(49),
    to_slogic(82),
    to_slogic(116),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(155),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(177),
    to_slogic(187),
    to_slogic(182),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(205),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(213),
    to_slogic(141),
    to_slogic(88),
    to_slogic(101),
    to_slogic(101),
    to_slogic(107),
    to_slogic(107),
    to_slogic(107),
    to_slogic(101),
    to_slogic(88),
    to_slogic(96),
    to_slogic(82),
    to_slogic(82),
    to_slogic(75),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(130),
    to_slogic(197),
    to_slogic(203),
    to_slogic(196),
    to_slogic(169),
    to_slogic(161),
    to_slogic(191),
    to_slogic(213),
    to_slogic(213),
    to_slogic(203),
    to_slogic(184),
    to_slogic(136),
    to_slogic(89),
    to_slogic(64),
    to_slogic(56),
    to_slogic(63),
    to_slogic(76),
    to_slogic(75),
    to_slogic(75),
    to_slogic(70),
    to_slogic(82),
    to_slogic(83),
    to_slogic(107),
    to_slogic(109),
    to_slogic(96),
    to_slogic(83),
    to_slogic(83),
    to_slogic(83),
    to_slogic(83),
    to_slogic(83),
    to_slogic(96),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(83),
    to_slogic(82),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(96),
    to_slogic(96),
    to_slogic(82),
    to_slogic(91),
    to_slogic(91),
    to_slogic(114),
    to_slogic(149),
    to_slogic(170),
    to_slogic(177),
    to_slogic(189),
    to_slogic(170),
    to_slogic(149),
    to_slogic(91),
    to_slogic(75),
    to_slogic(102),
    to_slogic(143),
    to_slogic(157),
    to_slogic(165),
    to_slogic(178),
    to_slogic(178),
    to_slogic(176),
    to_slogic(178),
    to_slogic(176),
    to_slogic(183),
    to_slogic(176),
    to_slogic(165),
    to_slogic(135),
    to_slogic(101),
    to_slogic(121),
    to_slogic(101),
    to_slogic(63),
    to_slogic(40),
    to_slogic(42),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(68),
    to_slogic(63),
    to_slogic(63),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(81),
    to_slogic(122),
    to_slogic(145),
    to_slogic(153),
    to_slogic(115),
    to_slogic(97),
    to_slogic(102),
    to_slogic(119),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(40),
    to_slogic(44),
    to_slogic(33),
    to_slogic(62),
    to_slogic(75),
    to_slogic(75),
    to_slogic(97),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(109),
    to_slogic(76),
    to_slogic(44),
    to_slogic(49),
    to_slogic(70),
    to_slogic(109),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(151),
    to_slogic(165),
    to_slogic(155),
    to_slogic(173),
    to_slogic(173),
    to_slogic(173),
    to_slogic(172),
    to_slogic(183),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(196),
    to_slogic(200),
    to_slogic(200),
    to_slogic(211),
    to_slogic(200),
    to_slogic(211),
    to_slogic(205),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(213),
    to_slogic(176),
    to_slogic(82),
    to_slogic(92),
    to_slogic(101),
    to_slogic(107),
    to_slogic(101),
    to_slogic(102),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(92),
    to_slogic(91),
    to_slogic(75),
    to_slogic(75),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(33),
    to_slogic(40),
    to_slogic(49),
    to_slogic(136),
    to_slogic(191),
    to_slogic(203),
    to_slogic(196),
    to_slogic(169),
    to_slogic(175),
    to_slogic(196),
    to_slogic(203),
    to_slogic(203),
    to_slogic(196),
    to_slogic(144),
    to_slogic(89),
    to_slogic(62),
    to_slogic(56),
    to_slogic(62),
    to_slogic(64),
    to_slogic(75),
    to_slogic(76),
    to_slogic(70),
    to_slogic(77),
    to_slogic(83),
    to_slogic(101),
    to_slogic(110),
    to_slogic(101),
    to_slogic(83),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(83),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(91),
    to_slogic(82),
    to_slogic(68),
    to_slogic(64),
    to_slogic(62),
    to_slogic(64),
    to_slogic(82),
    to_slogic(88),
    to_slogic(96),
    to_slogic(96),
    to_slogic(102),
    to_slogic(119),
    to_slogic(153),
    to_slogic(170),
    to_slogic(191),
    to_slogic(177),
    to_slogic(176),
    to_slogic(149),
    to_slogic(102),
    to_slogic(82),
    to_slogic(109),
    to_slogic(135),
    to_slogic(152),
    to_slogic(173),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(176),
    to_slogic(172),
    to_slogic(130),
    to_slogic(101),
    to_slogic(120),
    to_slogic(96),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(68),
    to_slogic(68),
    to_slogic(63),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(71),
    to_slogic(71),
    to_slogic(89),
    to_slogic(120),
    to_slogic(130),
    to_slogic(102),
    to_slogic(102),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(33),
    to_slogic(33),
    to_slogic(40),
    to_slogic(49),
    to_slogic(62),
    to_slogic(62),
    to_slogic(81),
    to_slogic(89),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(109),
    to_slogic(76),
    to_slogic(33),
    to_slogic(40),
    to_slogic(75),
    to_slogic(100),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(130),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(155),
    to_slogic(162),
    to_slogic(165),
    to_slogic(162),
    to_slogic(173),
    to_slogic(172),
    to_slogic(177),
    to_slogic(187),
    to_slogic(182),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(198),
    to_slogic(96),
    to_slogic(88),
    to_slogic(96),
    to_slogic(107),
    to_slogic(107),
    to_slogic(107),
    to_slogic(107),
    to_slogic(102),
    to_slogic(101),
    to_slogic(88),
    to_slogic(91),
    to_slogic(82),
    to_slogic(82),
    to_slogic(75),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(124),
    to_slogic(184),
    to_slogic(196),
    to_slogic(203),
    to_slogic(184),
    to_slogic(184),
    to_slogic(196),
    to_slogic(196),
    to_slogic(184),
    to_slogic(156),
    to_slogic(94),
    to_slogic(62),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(70),
    to_slogic(75),
    to_slogic(62),
    to_slogic(75),
    to_slogic(82),
    to_slogic(102),
    to_slogic(101),
    to_slogic(101),
    to_slogic(91),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(83),
    to_slogic(96),
    to_slogic(109),
    to_slogic(110),
    to_slogic(102),
    to_slogic(96),
    to_slogic(83),
    to_slogic(83),
    to_slogic(75),
    to_slogic(64),
    to_slogic(64),
    to_slogic(64),
    to_slogic(83),
    to_slogic(91),
    to_slogic(96),
    to_slogic(102),
    to_slogic(109),
    to_slogic(133),
    to_slogic(153),
    to_slogic(170),
    to_slogic(177),
    to_slogic(177),
    to_slogic(176),
    to_slogic(149),
    to_slogic(102),
    to_slogic(88),
    to_slogic(100),
    to_slogic(135),
    to_slogic(157),
    to_slogic(165),
    to_slogic(178),
    to_slogic(173),
    to_slogic(176),
    to_slogic(176),
    to_slogic(183),
    to_slogic(176),
    to_slogic(176),
    to_slogic(165),
    to_slogic(130),
    to_slogic(101),
    to_slogic(119),
    to_slogic(96),
    to_slogic(64),
    to_slogic(42),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(50),
    to_slogic(56),
    to_slogic(81),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(68),
    to_slogic(71),
    to_slogic(42),
    to_slogic(63),
    to_slogic(71),
    to_slogic(50),
    to_slogic(56),
    to_slogic(95),
    to_slogic(56),
    to_slogic(76),
    to_slogic(89),
    to_slogic(97),
    to_slogic(95),
    to_slogic(130),
    to_slogic(119),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(33),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(75),
    to_slogic(100),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(62),
    to_slogic(44),
    to_slogic(49),
    to_slogic(70),
    to_slogic(100),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(135),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(165),
    to_slogic(155),
    to_slogic(165),
    to_slogic(162),
    to_slogic(162),
    to_slogic(173),
    to_slogic(177),
    to_slogic(177),
    to_slogic(187),
    to_slogic(193),
    to_slogic(189),
    to_slogic(200),
    to_slogic(196),
    to_slogic(204),
    to_slogic(211),
    to_slogic(200),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(213),
    to_slogic(125),
    to_slogic(89),
    to_slogic(88),
    to_slogic(101),
    to_slogic(107),
    to_slogic(107),
    to_slogic(102),
    to_slogic(107),
    to_slogic(102),
    to_slogic(96),
    to_slogic(96),
    to_slogic(88),
    to_slogic(88),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(62),
    to_slogic(64),
    to_slogic(70),
    to_slogic(116),
    to_slogic(178),
    to_slogic(203),
    to_slogic(205),
    to_slogic(197),
    to_slogic(191),
    to_slogic(184),
    to_slogic(169),
    to_slogic(144),
    to_slogic(102),
    to_slogic(70),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(70),
    to_slogic(70),
    to_slogic(62),
    to_slogic(70),
    to_slogic(82),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(83),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(83),
    to_slogic(96),
    to_slogic(101),
    to_slogic(110),
    to_slogic(109),
    to_slogic(101),
    to_slogic(91),
    to_slogic(81),
    to_slogic(82),
    to_slogic(68),
    to_slogic(56),
    to_slogic(64),
    to_slogic(68),
    to_slogic(75),
    to_slogic(88),
    to_slogic(102),
    to_slogic(109),
    to_slogic(119),
    to_slogic(119),
    to_slogic(153),
    to_slogic(176),
    to_slogic(177),
    to_slogic(176),
    to_slogic(176),
    to_slogic(158),
    to_slogic(102),
    to_slogic(82),
    to_slogic(109),
    to_slogic(135),
    to_slogic(150),
    to_slogic(165),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(183),
    to_slogic(176),
    to_slogic(172),
    to_slogic(130),
    to_slogic(96),
    to_slogic(120),
    to_slogic(89),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(40),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(71),
    to_slogic(71),
    to_slogic(71),
    to_slogic(49),
    to_slogic(63),
    to_slogic(89),
    to_slogic(71),
    to_slogic(49),
    to_slogic(49),
    to_slogic(42),
    to_slogic(71),
    to_slogic(89),
    to_slogic(63),
    to_slogic(56),
    to_slogic(81),
    to_slogic(56),
    to_slogic(63),
    to_slogic(81),
    to_slogic(83),
    to_slogic(76),
    to_slogic(120),
    to_slogic(122),
    to_slogic(71),
    to_slogic(68),
    to_slogic(89),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(33),
    to_slogic(33),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(75),
    to_slogic(89),
    to_slogic(100),
    to_slogic(100),
    to_slogic(102),
    to_slogic(109),
    to_slogic(75),
    to_slogic(44),
    to_slogic(40),
    to_slogic(49),
    to_slogic(89),
    to_slogic(100),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(135),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(157),
    to_slogic(151),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(162),
    to_slogic(173),
    to_slogic(165),
    to_slogic(173),
    to_slogic(177),
    to_slogic(182),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(213),
    to_slogic(158),
    to_slogic(75),
    to_slogic(88),
    to_slogic(101),
    to_slogic(102),
    to_slogic(107),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(88),
    to_slogic(101),
    to_slogic(96),
    to_slogic(96),
    to_slogic(82),
    to_slogic(82),
    to_slogic(75),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(124),
    to_slogic(183),
    to_slogic(205),
    to_slogic(207),
    to_slogic(203),
    to_slogic(184),
    to_slogic(161),
    to_slogic(118),
    to_slogic(94),
    to_slogic(70),
    to_slogic(62),
    to_slogic(49),
    to_slogic(64),
    to_slogic(64),
    to_slogic(75),
    to_slogic(70),
    to_slogic(63),
    to_slogic(83),
    to_slogic(92),
    to_slogic(101),
    to_slogic(109),
    to_slogic(96),
    to_slogic(83),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(83),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(91),
    to_slogic(91),
    to_slogic(82),
    to_slogic(75),
    to_slogic(64),
    to_slogic(64),
    to_slogic(75),
    to_slogic(56),
    to_slogic(64),
    to_slogic(83),
    to_slogic(102),
    to_slogic(114),
    to_slogic(109),
    to_slogic(119),
    to_slogic(143),
    to_slogic(162),
    to_slogic(176),
    to_slogic(177),
    to_slogic(170),
    to_slogic(149),
    to_slogic(102),
    to_slogic(88),
    to_slogic(102),
    to_slogic(135),
    to_slogic(157),
    to_slogic(165),
    to_slogic(178),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(176),
    to_slogic(165),
    to_slogic(144),
    to_slogic(83),
    to_slogic(110),
    to_slogic(89),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(42),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(68),
    to_slogic(50),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(71),
    to_slogic(83),
    to_slogic(81),
    to_slogic(50),
    to_slogic(65),
    to_slogic(89),
    to_slogic(81),
    to_slogic(56),
    to_slogic(40),
    to_slogic(49),
    to_slogic(68),
    to_slogic(81),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(97),
    to_slogic(56),
    to_slogic(58),
    to_slogic(71),
    to_slogic(76),
    to_slogic(89),
    to_slogic(143),
    to_slogic(89),
    to_slogic(63),
    to_slogic(63),
    to_slogic(71),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(33),
    to_slogic(33),
    to_slogic(56),
    to_slogic(75),
    to_slogic(89),
    to_slogic(89),
    to_slogic(89),
    to_slogic(89),
    to_slogic(62),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(75),
    to_slogic(97),
    to_slogic(109),
    to_slogic(115),
    to_slogic(116),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(135),
    to_slogic(134),
    to_slogic(135),
    to_slogic(139),
    to_slogic(130),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(135),
    to_slogic(135),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(162),
    to_slogic(155),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(172),
    to_slogic(177),
    to_slogic(176),
    to_slogic(187),
    to_slogic(187),
    to_slogic(191),
    to_slogic(195),
    to_slogic(196),
    to_slogic(200),
    to_slogic(197),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(214),
    to_slogic(185),
    to_slogic(89),
    to_slogic(88),
    to_slogic(96),
    to_slogic(101),
    to_slogic(107),
    to_slogic(102),
    to_slogic(102),
    to_slogic(101),
    to_slogic(96),
    to_slogic(101),
    to_slogic(96),
    to_slogic(91),
    to_slogic(83),
    to_slogic(96),
    to_slogic(91),
    to_slogic(83),
    to_slogic(94),
    to_slogic(92),
    to_slogic(126),
    to_slogic(177),
    to_slogic(205),
    to_slogic(207),
    to_slogic(196),
    to_slogic(161),
    to_slogic(107),
    to_slogic(89),
    to_slogic(70),
    to_slogic(64),
    to_slogic(62),
    to_slogic(63),
    to_slogic(75),
    to_slogic(75),
    to_slogic(70),
    to_slogic(70),
    to_slogic(82),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(101),
    to_slogic(91),
    to_slogic(75),
    to_slogic(70),
    to_slogic(69),
    to_slogic(75),
    to_slogic(88),
    to_slogic(91),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(101),
    to_slogic(101),
    to_slogic(91),
    to_slogic(82),
    to_slogic(64),
    to_slogic(64),
    to_slogic(64),
    to_slogic(68),
    to_slogic(64),
    to_slogic(40),
    to_slogic(82),
    to_slogic(96),
    to_slogic(96),
    to_slogic(102),
    to_slogic(114),
    to_slogic(143),
    to_slogic(165),
    to_slogic(177),
    to_slogic(177),
    to_slogic(176),
    to_slogic(149),
    to_slogic(118),
    to_slogic(88),
    to_slogic(109),
    to_slogic(130),
    to_slogic(152),
    to_slogic(165),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(172),
    to_slogic(172),
    to_slogic(144),
    to_slogic(87),
    to_slogic(101),
    to_slogic(83),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(81),
    to_slogic(81),
    to_slogic(89),
    to_slogic(49),
    to_slogic(71),
    to_slogic(95),
    to_slogic(89),
    to_slogic(81),
    to_slogic(42),
    to_slogic(50),
    to_slogic(49),
    to_slogic(95),
    to_slogic(50),
    to_slogic(49),
    to_slogic(63),
    to_slogic(113),
    to_slogic(71),
    to_slogic(63),
    to_slogic(58),
    to_slogic(84),
    to_slogic(97),
    to_slogic(138),
    to_slogic(127),
    to_slogic(71),
    to_slogic(63),
    to_slogic(68),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(62),
    to_slogic(62),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(62),
    to_slogic(76),
    to_slogic(89),
    to_slogic(100),
    to_slogic(100),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(135),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(165),
    to_slogic(157),
    to_slogic(173),
    to_slogic(165),
    to_slogic(178),
    to_slogic(172),
    to_slogic(177),
    to_slogic(182),
    to_slogic(182),
    to_slogic(193),
    to_slogic(195),
    to_slogic(196),
    to_slogic(200),
    to_slogic(211),
    to_slogic(205),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(213),
    to_slogic(204),
    to_slogic(107),
    to_slogic(82),
    to_slogic(88),
    to_slogic(88),
    to_slogic(101),
    to_slogic(101),
    to_slogic(107),
    to_slogic(107),
    to_slogic(101),
    to_slogic(102),
    to_slogic(101),
    to_slogic(101),
    to_slogic(91),
    to_slogic(96),
    to_slogic(101),
    to_slogic(101),
    to_slogic(94),
    to_slogic(96),
    to_slogic(118),
    to_slogic(165),
    to_slogic(191),
    to_slogic(191),
    to_slogic(161),
    to_slogic(116),
    to_slogic(88),
    to_slogic(82),
    to_slogic(82),
    to_slogic(64),
    to_slogic(70),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(87),
    to_slogic(107),
    to_slogic(109),
    to_slogic(109),
    to_slogic(83),
    to_slogic(82),
    to_slogic(82),
    to_slogic(64),
    to_slogic(64),
    to_slogic(75),
    to_slogic(96),
    to_slogic(101),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(102),
    to_slogic(96),
    to_slogic(88),
    to_slogic(64),
    to_slogic(64),
    to_slogic(75),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(49),
    to_slogic(64),
    to_slogic(82),
    to_slogic(91),
    to_slogic(89),
    to_slogic(102),
    to_slogic(133),
    to_slogic(162),
    to_slogic(176),
    to_slogic(177),
    to_slogic(170),
    to_slogic(158),
    to_slogic(119),
    to_slogic(88),
    to_slogic(109),
    to_slogic(130),
    to_slogic(151),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(183),
    to_slogic(183),
    to_slogic(178),
    to_slogic(165),
    to_slogic(152),
    to_slogic(83),
    to_slogic(87),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(81),
    to_slogic(50),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(81),
    to_slogic(71),
    to_slogic(42),
    to_slogic(71),
    to_slogic(97),
    to_slogic(115),
    to_slogic(102),
    to_slogic(68),
    to_slogic(56),
    to_slogic(50),
    to_slogic(81),
    to_slogic(71),
    to_slogic(49),
    to_slogic(56),
    to_slogic(68),
    to_slogic(115),
    to_slogic(71),
    to_slogic(56),
    to_slogic(76),
    to_slogic(109),
    to_slogic(115),
    to_slogic(152),
    to_slogic(107),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(64),
    to_slogic(89),
    to_slogic(92),
    to_slogic(102),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(134),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(143),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(173),
    to_slogic(172),
    to_slogic(177),
    to_slogic(176),
    to_slogic(182),
    to_slogic(187),
    to_slogic(189),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(205),
    to_slogic(211),
    to_slogic(208),
    to_slogic(211),
    to_slogic(208),
    to_slogic(214),
    to_slogic(214),
    to_slogic(207),
    to_slogic(133),
    to_slogic(82),
    to_slogic(82),
    to_slogic(94),
    to_slogic(96),
    to_slogic(102),
    to_slogic(101),
    to_slogic(102),
    to_slogic(107),
    to_slogic(107),
    to_slogic(102),
    to_slogic(101),
    to_slogic(96),
    to_slogic(107),
    to_slogic(107),
    to_slogic(107),
    to_slogic(107),
    to_slogic(109),
    to_slogic(109),
    to_slogic(136),
    to_slogic(144),
    to_slogic(143),
    to_slogic(102),
    to_slogic(88),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(89),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(83),
    to_slogic(101),
    to_slogic(109),
    to_slogic(107),
    to_slogic(88),
    to_slogic(75),
    to_slogic(75),
    to_slogic(64),
    to_slogic(63),
    to_slogic(75),
    to_slogic(83),
    to_slogic(101),
    to_slogic(109),
    to_slogic(120),
    to_slogic(114),
    to_slogic(109),
    to_slogic(101),
    to_slogic(91),
    to_slogic(68),
    to_slogic(64),
    to_slogic(64),
    to_slogic(64),
    to_slogic(64),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(83),
    to_slogic(83),
    to_slogic(102),
    to_slogic(119),
    to_slogic(153),
    to_slogic(170),
    to_slogic(176),
    to_slogic(176),
    to_slogic(153),
    to_slogic(130),
    to_slogic(101),
    to_slogic(102),
    to_slogic(130),
    to_slogic(152),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(165),
    to_slogic(157),
    to_slogic(92),
    to_slogic(68),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(83),
    to_slogic(63),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(65),
    to_slogic(89),
    to_slogic(63),
    to_slogic(42),
    to_slogic(58),
    to_slogic(97),
    to_slogic(113),
    to_slogic(107),
    to_slogic(71),
    to_slogic(42),
    to_slogic(56),
    to_slogic(71),
    to_slogic(113),
    to_slogic(49),
    to_slogic(36),
    to_slogic(65),
    to_slogic(89),
    to_slogic(89),
    to_slogic(65),
    to_slogic(65),
    to_slogic(115),
    to_slogic(115),
    to_slogic(95),
    to_slogic(113),
    to_slogic(97),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(62),
    to_slogic(62),
    to_slogic(75),
    to_slogic(89),
    to_slogic(97),
    to_slogic(97),
    to_slogic(109),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(143),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(162),
    to_slogic(162),
    to_slogic(165),
    to_slogic(177),
    to_slogic(177),
    to_slogic(182),
    to_slogic(187),
    to_slogic(187),
    to_slogic(189),
    to_slogic(193),
    to_slogic(200),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(211),
    to_slogic(214),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(213),
    to_slogic(167),
    to_slogic(82),
    to_slogic(82),
    to_slogic(91),
    to_slogic(88),
    to_slogic(96),
    to_slogic(101),
    to_slogic(107),
    to_slogic(107),
    to_slogic(102),
    to_slogic(109),
    to_slogic(102),
    to_slogic(107),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(107),
    to_slogic(107),
    to_slogic(101),
    to_slogic(116),
    to_slogic(118),
    to_slogic(107),
    to_slogic(96),
    to_slogic(82),
    to_slogic(92),
    to_slogic(82),
    to_slogic(92),
    to_slogic(92),
    to_slogic(82),
    to_slogic(89),
    to_slogic(70),
    to_slogic(75),
    to_slogic(82),
    to_slogic(96),
    to_slogic(109),
    to_slogic(96),
    to_slogic(91),
    to_slogic(82),
    to_slogic(75),
    to_slogic(64),
    to_slogic(64),
    to_slogic(64),
    to_slogic(75),
    to_slogic(101),
    to_slogic(109),
    to_slogic(110),
    to_slogic(120),
    to_slogic(120),
    to_slogic(102),
    to_slogic(96),
    to_slogic(91),
    to_slogic(75),
    to_slogic(64),
    to_slogic(64),
    to_slogic(62),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(91),
    to_slogic(81),
    to_slogic(119),
    to_slogic(153),
    to_slogic(176),
    to_slogic(177),
    to_slogic(176),
    to_slogic(158),
    to_slogic(130),
    to_slogic(102),
    to_slogic(107),
    to_slogic(130),
    to_slogic(151),
    to_slogic(158),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(165),
    to_slogic(157),
    to_slogic(83),
    to_slogic(69),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(68),
    to_slogic(81),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(68),
    to_slogic(95),
    to_slogic(56),
    to_slogic(42),
    to_slogic(56),
    to_slogic(97),
    to_slogic(89),
    to_slogic(120),
    to_slogic(89),
    to_slogic(42),
    to_slogic(42),
    to_slogic(83),
    to_slogic(113),
    to_slogic(89),
    to_slogic(36),
    to_slogic(56),
    to_slogic(71),
    to_slogic(102),
    to_slogic(63),
    to_slogic(71),
    to_slogic(97),
    to_slogic(107),
    to_slogic(107),
    to_slogic(83),
    to_slogic(95),
    to_slogic(68),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(40),
    to_slogic(33),
    to_slogic(33),
    to_slogic(44),
    to_slogic(56),
    to_slogic(62),
    to_slogic(62),
    to_slogic(89),
    to_slogic(89),
    to_slogic(100),
    to_slogic(109),
    to_slogic(97),
    to_slogic(121),
    to_slogic(109),
    to_slogic(121),
    to_slogic(126),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(135),
    to_slogic(130),
    to_slogic(139),
    to_slogic(139),
    to_slogic(143),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(135),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(155),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(172),
    to_slogic(172),
    to_slogic(183),
    to_slogic(182),
    to_slogic(187),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(214),
    to_slogic(214),
    to_slogic(189),
    to_slogic(96),
    to_slogic(82),
    to_slogic(88),
    to_slogic(91),
    to_slogic(96),
    to_slogic(102),
    to_slogic(102),
    to_slogic(107),
    to_slogic(118),
    to_slogic(102),
    to_slogic(109),
    to_slogic(107),
    to_slogic(118),
    to_slogic(118),
    to_slogic(118),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(96),
    to_slogic(96),
    to_slogic(92),
    to_slogic(96),
    to_slogic(96),
    to_slogic(94),
    to_slogic(96),
    to_slogic(82),
    to_slogic(81),
    to_slogic(82),
    to_slogic(82),
    to_slogic(87),
    to_slogic(109),
    to_slogic(96),
    to_slogic(91),
    to_slogic(82),
    to_slogic(82),
    to_slogic(75),
    to_slogic(64),
    to_slogic(64),
    to_slogic(75),
    to_slogic(91),
    to_slogic(109),
    to_slogic(109),
    to_slogic(120),
    to_slogic(119),
    to_slogic(109),
    to_slogic(101),
    to_slogic(96),
    to_slogic(82),
    to_slogic(64),
    to_slogic(64),
    to_slogic(56),
    to_slogic(64),
    to_slogic(62),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(64),
    to_slogic(64),
    to_slogic(64),
    to_slogic(68),
    to_slogic(81),
    to_slogic(114),
    to_slogic(153),
    to_slogic(177),
    to_slogic(196),
    to_slogic(196),
    to_slogic(176),
    to_slogic(143),
    to_slogic(102),
    to_slogic(109),
    to_slogic(130),
    to_slogic(151),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(183),
    to_slogic(178),
    to_slogic(165),
    to_slogic(118),
    to_slogic(69),
    to_slogic(56),
    to_slogic(68),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(89),
    to_slogic(56),
    to_slogic(42),
    to_slogic(42),
    to_slogic(71),
    to_slogic(89),
    to_slogic(42),
    to_slogic(42),
    to_slogic(50),
    to_slogic(102),
    to_slogic(84),
    to_slogic(102),
    to_slogic(127),
    to_slogic(56),
    to_slogic(42),
    to_slogic(63),
    to_slogic(102),
    to_slogic(113),
    to_slogic(56),
    to_slogic(36),
    to_slogic(63),
    to_slogic(89),
    to_slogic(102),
    to_slogic(50),
    to_slogic(71),
    to_slogic(102),
    to_slogic(115),
    to_slogic(95),
    to_slogic(68),
    to_slogic(63),
    to_slogic(40),
    to_slogic(40),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(44),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(89),
    to_slogic(97),
    to_slogic(97),
    to_slogic(109),
    to_slogic(109),
    to_slogic(121),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(134),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(162),
    to_slogic(173),
    to_slogic(172),
    to_slogic(177),
    to_slogic(176),
    to_slogic(182),
    to_slogic(187),
    to_slogic(185),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(213),
    to_slogic(207),
    to_slogic(109),
    to_slogic(64),
    to_slogic(88),
    to_slogic(88),
    to_slogic(101),
    to_slogic(102),
    to_slogic(107),
    to_slogic(109),
    to_slogic(118),
    to_slogic(109),
    to_slogic(120),
    to_slogic(118),
    to_slogic(118),
    to_slogic(118),
    to_slogic(116),
    to_slogic(107),
    to_slogic(116),
    to_slogic(109),
    to_slogic(102),
    to_slogic(101),
    to_slogic(100),
    to_slogic(100),
    to_slogic(94),
    to_slogic(101),
    to_slogic(116),
    to_slogic(109),
    to_slogic(99),
    to_slogic(82),
    to_slogic(82),
    to_slogic(82),
    to_slogic(96),
    to_slogic(91),
    to_slogic(91),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(101),
    to_slogic(109),
    to_slogic(114),
    to_slogic(120),
    to_slogic(114),
    to_slogic(102),
    to_slogic(96),
    to_slogic(88),
    to_slogic(64),
    to_slogic(64),
    to_slogic(62),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(68),
    to_slogic(114),
    to_slogic(165),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(193),
    to_slogic(171),
    to_slogic(118),
    to_slogic(107),
    to_slogic(135),
    to_slogic(152),
    to_slogic(165),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(183),
    to_slogic(183),
    to_slogic(178),
    to_slogic(157),
    to_slogic(101),
    to_slogic(69),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(42),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(50),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(50),
    to_slogic(71),
    to_slogic(71),
    to_slogic(42),
    to_slogic(50),
    to_slogic(95),
    to_slogic(102),
    to_slogic(50),
    to_slogic(50),
    to_slogic(50),
    to_slogic(102),
    to_slogic(91),
    to_slogic(75),
    to_slogic(130),
    to_slogic(97),
    to_slogic(56),
    to_slogic(50),
    to_slogic(95),
    to_slogic(102),
    to_slogic(71),
    to_slogic(40),
    to_slogic(42),
    to_slogic(71),
    to_slogic(114),
    to_slogic(83),
    to_slogic(42),
    to_slogic(71),
    to_slogic(97),
    to_slogic(107),
    to_slogic(65),
    to_slogic(56),
    to_slogic(49),
    to_slogic(33),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(62),
    to_slogic(89),
    to_slogic(97),
    to_slogic(97),
    to_slogic(109),
    to_slogic(109),
    to_slogic(121),
    to_slogic(109),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(135),
    to_slogic(121),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(146),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(151),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(162),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(177),
    to_slogic(176),
    to_slogic(183),
    to_slogic(182),
    to_slogic(182),
    to_slogic(187),
    to_slogic(191),
    to_slogic(200),
    to_slogic(196),
    to_slogic(200),
    to_slogic(211),
    to_slogic(205),
    to_slogic(211),
    to_slogic(211),
    to_slogic(205),
    to_slogic(214),
    to_slogic(211),
    to_slogic(132),
    to_slogic(82),
    to_slogic(82),
    to_slogic(88),
    to_slogic(91),
    to_slogic(101),
    to_slogic(102),
    to_slogic(107),
    to_slogic(107),
    to_slogic(118),
    to_slogic(118),
    to_slogic(118),
    to_slogic(128),
    to_slogic(118),
    to_slogic(116),
    to_slogic(116),
    to_slogic(118),
    to_slogic(107),
    to_slogic(116),
    to_slogic(109),
    to_slogic(101),
    to_slogic(101),
    to_slogic(109),
    to_slogic(116),
    to_slogic(107),
    to_slogic(102),
    to_slogic(96),
    to_slogic(92),
    to_slogic(82),
    to_slogic(96),
    to_slogic(96),
    to_slogic(101),
    to_slogic(91),
    to_slogic(82),
    to_slogic(64),
    to_slogic(75),
    to_slogic(64),
    to_slogic(75),
    to_slogic(75),
    to_slogic(83),
    to_slogic(96),
    to_slogic(109),
    to_slogic(120),
    to_slogic(125),
    to_slogic(121),
    to_slogic(109),
    to_slogic(102),
    to_slogic(91),
    to_slogic(82),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(64),
    to_slogic(63),
    to_slogic(119),
    to_slogic(177),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(193),
    to_slogic(176),
    to_slogic(125),
    to_slogic(107),
    to_slogic(126),
    to_slogic(151),
    to_slogic(165),
    to_slogic(173),
    to_slogic(176),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(158),
    to_slogic(134),
    to_slogic(96),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(49),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(89),
    to_slogic(42),
    to_slogic(42),
    to_slogic(113),
    to_slogic(89),
    to_slogic(50),
    to_slogic(50),
    to_slogic(56),
    to_slogic(107),
    to_slogic(84),
    to_slogic(76),
    to_slogic(127),
    to_slogic(120),
    to_slogic(56),
    to_slogic(42),
    to_slogic(56),
    to_slogic(102),
    to_slogic(63),
    to_slogic(63),
    to_slogic(42),
    to_slogic(69),
    to_slogic(81),
    to_slogic(107),
    to_slogic(50),
    to_slogic(71),
    to_slogic(75),
    to_slogic(107),
    to_slogic(89),
    to_slogic(89),
    to_slogic(56),
    to_slogic(40),
    to_slogic(33),
    to_slogic(33),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(81),
    to_slogic(97),
    to_slogic(97),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(135),
    to_slogic(135),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(157),
    to_slogic(165),
    to_slogic(165),
    to_slogic(173),
    to_slogic(165),
    to_slogic(172),
    to_slogic(177),
    to_slogic(177),
    to_slogic(177),
    to_slogic(187),
    to_slogic(189),
    to_slogic(193),
    to_slogic(195),
    to_slogic(200),
    to_slogic(200),
    to_slogic(205),
    to_slogic(200),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(213),
    to_slogic(165),
    to_slogic(75),
    to_slogic(75),
    to_slogic(88),
    to_slogic(96),
    to_slogic(101),
    to_slogic(102),
    to_slogic(102),
    to_slogic(109),
    to_slogic(109),
    to_slogic(118),
    to_slogic(118),
    to_slogic(118),
    to_slogic(116),
    to_slogic(118),
    to_slogic(116),
    to_slogic(116),
    to_slogic(116),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(116),
    to_slogic(116),
    to_slogic(121),
    to_slogic(116),
    to_slogic(109),
    to_slogic(99),
    to_slogic(96),
    to_slogic(96),
    to_slogic(96),
    to_slogic(96),
    to_slogic(91),
    to_slogic(83),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(82),
    to_slogic(75),
    to_slogic(82),
    to_slogic(96),
    to_slogic(109),
    to_slogic(120),
    to_slogic(126),
    to_slogic(119),
    to_slogic(109),
    to_slogic(102),
    to_slogic(91),
    to_slogic(82),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(62),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(64),
    to_slogic(82),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(119),
    to_slogic(185),
    to_slogic(196),
    to_slogic(204),
    to_slogic(204),
    to_slogic(193),
    to_slogic(189),
    to_slogic(144),
    to_slogic(107),
    to_slogic(130),
    to_slogic(152),
    to_slogic(165),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(183),
    to_slogic(173),
    to_slogic(165),
    to_slogic(127),
    to_slogic(96),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(56),
    to_slogic(56),
    to_slogic(75),
    to_slogic(75),
    to_slogic(68),
    to_slogic(50),
    to_slogic(75),
    to_slogic(63),
    to_slogic(50),
    to_slogic(120),
    to_slogic(75),
    to_slogic(56),
    to_slogic(50),
    to_slogic(65),
    to_slogic(107),
    to_slogic(83),
    to_slogic(76),
    to_slogic(81),
    to_slogic(138),
    to_slogic(83),
    to_slogic(42),
    to_slogic(56),
    to_slogic(102),
    to_slogic(97),
    to_slogic(56),
    to_slogic(63),
    to_slogic(63),
    to_slogic(81),
    to_slogic(68),
    to_slogic(71),
    to_slogic(56),
    to_slogic(71),
    to_slogic(107),
    to_slogic(84),
    to_slogic(115),
    to_slogic(95),
    to_slogic(49),
    to_slogic(33),
    to_slogic(44),
    to_slogic(44),
    to_slogic(62),
    to_slogic(81),
    to_slogic(89),
    to_slogic(97),
    to_slogic(97),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(121),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(121),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(134),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(144),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(146),
    to_slogic(151),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(151),
    to_slogic(157),
    to_slogic(165),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(173),
    to_slogic(177),
    to_slogic(177),
    to_slogic(182),
    to_slogic(187),
    to_slogic(182),
    to_slogic(189),
    to_slogic(193),
    to_slogic(200),
    to_slogic(196),
    to_slogic(204),
    to_slogic(211),
    to_slogic(205),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(189),
    to_slogic(91),
    to_slogic(82),
    to_slogic(88),
    to_slogic(88),
    to_slogic(101),
    to_slogic(101),
    to_slogic(96),
    to_slogic(107),
    to_slogic(118),
    to_slogic(118),
    to_slogic(109),
    to_slogic(118),
    to_slogic(118),
    to_slogic(126),
    to_slogic(121),
    to_slogic(116),
    to_slogic(116),
    to_slogic(118),
    to_slogic(116),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(118),
    to_slogic(116),
    to_slogic(100),
    to_slogic(96),
    to_slogic(83),
    to_slogic(101),
    to_slogic(91),
    to_slogic(87),
    to_slogic(82),
    to_slogic(83),
    to_slogic(91),
    to_slogic(83),
    to_slogic(82),
    to_slogic(75),
    to_slogic(82),
    to_slogic(87),
    to_slogic(110),
    to_slogic(120),
    to_slogic(125),
    to_slogic(125),
    to_slogic(120),
    to_slogic(109),
    to_slogic(89),
    to_slogic(82),
    to_slogic(75),
    to_slogic(64),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(62),
    to_slogic(64),
    to_slogic(70),
    to_slogic(89),
    to_slogic(92),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(102),
    to_slogic(177),
    to_slogic(196),
    to_slogic(204),
    to_slogic(196),
    to_slogic(193),
    to_slogic(182),
    to_slogic(130),
    to_slogic(117),
    to_slogic(130),
    to_slogic(151),
    to_slogic(165),
    to_slogic(173),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(157),
    to_slogic(96),
    to_slogic(75),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(40),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(56),
    to_slogic(63),
    to_slogic(64),
    to_slogic(63),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(56),
    to_slogic(56),
    to_slogic(75),
    to_slogic(71),
    to_slogic(127),
    to_slogic(64),
    to_slogic(56),
    to_slogic(56),
    to_slogic(65),
    to_slogic(113),
    to_slogic(71),
    to_slogic(71),
    to_slogic(76),
    to_slogic(102),
    to_slogic(115),
    to_slogic(65),
    to_slogic(50),
    to_slogic(113),
    to_slogic(113),
    to_slogic(49),
    to_slogic(42),
    to_slogic(56),
    to_slogic(81),
    to_slogic(75),
    to_slogic(63),
    to_slogic(50),
    to_slogic(56),
    to_slogic(71),
    to_slogic(84),
    to_slogic(89),
    to_slogic(119),
    to_slogic(95),
    to_slogic(49),
    to_slogic(49),
    to_slogic(76),
    to_slogic(81),
    to_slogic(81),
    to_slogic(89),
    to_slogic(97),
    to_slogic(109),
    to_slogic(109),
    to_slogic(115),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(130),
    to_slogic(135),
    to_slogic(135),
    to_slogic(135),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(157),
    to_slogic(152),
    to_slogic(157),
    to_slogic(151),
    to_slogic(165),
    to_slogic(162),
    to_slogic(162),
    to_slogic(173),
    to_slogic(165),
    to_slogic(172),
    to_slogic(177),
    to_slogic(177),
    to_slogic(182),
    to_slogic(187),
    to_slogic(193),
    to_slogic(191),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(200),
    to_slogic(205),
    to_slogic(211),
    to_slogic(205),
    to_slogic(211),
    to_slogic(213),
    to_slogic(204),
    to_slogic(120),
    to_slogic(83),
    to_slogic(88),
    to_slogic(88),
    to_slogic(88),
    to_slogic(88),
    to_slogic(101),
    to_slogic(102),
    to_slogic(109),
    to_slogic(118),
    to_slogic(118),
    to_slogic(128),
    to_slogic(130),
    to_slogic(130),
    to_slogic(118),
    to_slogic(121),
    to_slogic(116),
    to_slogic(121),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(109),
    to_slogic(94),
    to_slogic(96),
    to_slogic(92),
    to_slogic(83),
    to_slogic(83),
    to_slogic(83),
    to_slogic(83),
    to_slogic(83),
    to_slogic(83),
    to_slogic(83),
    to_slogic(82),
    to_slogic(82),
    to_slogic(83),
    to_slogic(101),
    to_slogic(120),
    to_slogic(125),
    to_slogic(132),
    to_slogic(126),
    to_slogic(114),
    to_slogic(96),
    to_slogic(88),
    to_slogic(75),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(82),
    to_slogic(96),
    to_slogic(100),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(49),
    to_slogic(56),
    to_slogic(101),
    to_slogic(176),
    to_slogic(196),
    to_slogic(196),
    to_slogic(204),
    to_slogic(193),
    to_slogic(176),
    to_slogic(130),
    to_slogic(107),
    to_slogic(135),
    to_slogic(152),
    to_slogic(165),
    to_slogic(172),
    to_slogic(178),
    to_slogic(178),
    to_slogic(178),
    to_slogic(183),
    to_slogic(178),
    to_slogic(178),
    to_slogic(158),
    to_slogic(91),
    to_slogic(83),
    to_slogic(56),
    to_slogic(56),
    to_slogic(40),
    to_slogic(40),
    to_slogic(63),
    to_slogic(49),
    to_slogic(56),
    to_slogic(50),
    to_slogic(68),
    to_slogic(75),
    to_slogic(64),
    to_slogic(68),
    to_slogic(63),
    to_slogic(75),
    to_slogic(63),
    to_slogic(56),
    to_slogic(91),
    to_slogic(102),
    to_slogic(113),
    to_slogic(56),
    to_slogic(65),
    to_slogic(49),
    to_slogic(64),
    to_slogic(107),
    to_slogic(75),
    to_slogic(56),
    to_slogic(75),
    to_slogic(71),
    to_slogic(107),
    to_slogic(107),
    to_slogic(56),
    to_slogic(115),
    to_slogic(95),
    to_slogic(49),
    to_slogic(50),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(68),
    to_slogic(56),
    to_slogic(50),
    to_slogic(63),
    to_slogic(97),
    to_slogic(49),
    to_slogic(89),
    to_slogic(91),
    to_slogic(88),
    to_slogic(62),
    to_slogic(81),
    to_slogic(81),
    to_slogic(89),
    to_slogic(89),
    to_slogic(100),
    to_slogic(100),
    to_slogic(109),
    to_slogic(115),
    to_slogic(109),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(121),
    to_slogic(130),
    to_slogic(126),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(121),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(139),
    to_slogic(135),
    to_slogic(130),
    to_slogic(130),
    to_slogic(135),
    to_slogic(134),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(139),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(144),
    to_slogic(152),
    to_slogic(152),
    to_slogic(152),
    to_slogic(157),
    to_slogic(155),
    to_slogic(157),
    to_slogic(152),
    to_slogic(155),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(162),
    to_slogic(172),
    to_slogic(172),
    to_slogic(172),
    to_slogic(176),
    to_slogic(187),
    to_slogic(182),
    to_slogic(193),
    to_slogic(193),
    to_slogic(193),
    to_slogic(200),
    to_slogic(196),
    to_slogic(200),
    to_slogic(204),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(211),
    to_slogic(144),
    to_slogic(102),
    to_slogic(96),
    to_slogic(91),
    to_slogic(88),
    to_slogic(96),
    to_slogic(96),
    to_slogic(107),
    to_slogic(107),
    to_slogic(107),
    to_slogic(124),
    to_slogic(130),
    to_slogic(130),
    to_slogic(130),
    to_slogic(126),
    to_slogic(126),
    to_slogic(126),
    to_slogic(121),
    to_slogic(130),
    to_slogic(143),
    to_slogic(135),
    to_slogic(130),
    to_slogic(116),
    to_slogic(102),
    to_slogic(92),
    to_slogic(92),
    to_slogic(82),
    to_slogic(75),
    to_slogic(75),
    to_slogic(75),
    to_slogic(87),
    to_slogic(91),
    to_slogic(91),
    to_slogic(87),
    to_slogic(83),
    to_slogic(82),
    to_slogic(91),
    to_slogic(101),
    to_slogic(125),
    to_slogic(125),
    to_slogic(133),
    to_slogic(120),
    to_slogic(109),
    to_slogic(91),
    to_slogic(75),
    to_slogic(56),
    to_slogic(56),
    to_slogic(49),
    to_slogic(44),
    to_slogic(49),
    to_slogic(56),
    to_slogic(75),
    to_slogic(83),
    to_slogic(96),
    to_slogic(100),
    to_slogic(102)
  );
end package;
