library ieee;
use ieee.std_logic_1164.all;

library work;
use work.slogic_pkg.all;
use work.sobel_pkg.all;
